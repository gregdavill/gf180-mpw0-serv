* NGSPICE file created from serv_1.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__sdffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__sdffq_1 D SE SI CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_4 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyd_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyd_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnq_1 D CLKN Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_2 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_2 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

.subckt serv_1 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_oeb[0] io_oeb[1] io_oeb[2]
+ io_oeb[3] io_oeb[4] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] vdd vss
XFILLER_67_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05903_ _01528_ _01529_ _01530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__10669__A1 _05137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09671_ _04395_ _04396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06883_ u_cpu.rf_ram.memory\[116\]\[7\] u_cpu.rf_ram.memory\[117\]\[7\] u_cpu.rf_ram.memory\[118\]\[7\]
+ u_cpu.rf_ram.memory\[119\]\[7\] _02136_ _01707_ _02493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_80_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06337__A2 _01952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12595__CLK net274 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07534__A1 _02987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05834_ u_cpu.cpu.ctrl.o_ibus_adr\[7\] u_cpu.cpu.ctrl.o_ibus_adr\[6\] u_cpu.cpu.ctrl.o_ibus_adr\[5\]
+ _01464_ _01475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_08622_ _03285_ _02921_ _03711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09812__B _04531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout56_I net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05765_ u_cpu.cpu.immdec.imm24_20\[1\] _01388_ _01415_ _01416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08553_ _03484_ _03666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09287__A1 u_cpu.rf_ram.memory\[117\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11094__A1 _02684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07504_ _02987_ _02984_ _02988_ _00123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11094__B2 _01386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08484_ _03595_ _03621_ _03626_ _00465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_u_scanchain_local.scan_flop\[45\]_SE net559 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07837__A2 _03205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06896__I0 u_cpu.rf_ram.memory\[64\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10841__A1 _05209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07435_ _02889_ _02942_ _02944_ _00098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07366_ _02731_ _02891_ _02892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06317_ _01929_ _01931_ _01932_ _01933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09105_ _03969_ _04015_ _04017_ _00695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10185__S _04849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08262__A2 _03474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07297_ _02768_ _02834_ _02841_ _00063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09036_ _03971_ _03973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06248_ u_cpu.rf_ram.memory\[52\]\[1\] u_cpu.rf_ram.memory\[53\]\[1\] u_cpu.rf_ram.memory\[54\]\[1\]
+ u_cpu.rf_ram.memory\[55\]\[1\] _01863_ _01653_ _01864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_11_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08014__A2 _03324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06179_ _01791_ _01794_ _01795_ _01796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_2_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06415__I3 u_cpu.rf_ram.memory\[91\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06576__A2 _02188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11812__CLK net376 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09938_ _04578_ _04639_ _04423_ _04640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_63_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05806__I _01452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09869_ _04575_ _04580_ _04581_ _04583_ _04584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_3202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06328__A2 _01943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11900_ _00596_ net468 u_cpu.rf_ram.memory\[132\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11831_ _00527_ net478 u_cpu.rf_ram.memory\[138\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09278__A1 u_cpu.rf_ram.memory\[117\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11085__A1 _04026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11762_ _00458_ net490 u_cpu.rf_ram.memory\[141\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07828__A2 _03208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06187__S1 _01803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09013__I _03957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05839__A1 _01473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10713_ u_cpu.rf_ram.memory\[104\]\[4\] _05180_ _05183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11693_ _00397_ net331 u_cpu.rf_ram.memory\[56\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06500__A2 _02108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06351__I2 u_cpu.rf_ram.memory\[22\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10644_ _05137_ _05132_ _05139_ _01113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10575_ _03112_ _05097_ _01086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08253__A2 _03473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10060__A2 _04429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12314_ _00994_ net528 u_cpu.cpu.ctrl.o_ibus_adr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[34\] u_arbiter.i_wb_cpu_rdt\[31\] net549 u_arbiter.i_wb_cpu_dbus_dat\[28\]
+ net16 u_scanchain_local.module_data_in\[34\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__09202__A1 _02551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08005__A2 _03313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12245_ _00928_ net272 u_cpu.rf_ram.memory\[32\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10348__B1 _04945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12176_ _00859_ net387 u_arbiter.i_wb_cpu_dbus_dat\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10899__A1 _05300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06567__A2 _02179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11492__CLK net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08299__I _02776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11127_ _05445_ _05447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_46_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11058_ _05359_ _05392_ _05399_ _01267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_49_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11312__A2 _05558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10009_ u_cpu.cpu.immdec.imm30_25\[4\] _04667_ _04695_ u_cpu.cpu.immdec.imm30_25\[5\]
+ _04705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_36_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[68\]_SE net559 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout260_I net261 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout358_I net359 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11076__A1 _05357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10823__A1 _05211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout525_I net527 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08492__A2 _03622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07220_ u_cpu.rf_ram.memory\[21\]\[0\] _02793_ _02794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06893__I3 u_cpu.rf_ram.memory\[87\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07151_ _02732_ _02733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09441__A1 _04152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08244__A2 _03462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06102_ _01715_ _01718_ _01719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10051__A2 _04738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07082_ u_cpu.cpu.state.o_cnt_r\[0\] u_cpu.cpu.state.o_cnt_r\[1\] u_cpu.cpu.state.o_cnt_r\[2\]
+ _02563_ _02674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_69_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09992__A2 _04452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06033_ _01581_ _01650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout105 net107 net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout116 net119 net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__07755__A1 _03075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout127 net129 net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout138 net139 net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__10532__I _05071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout149 net151 net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_07984_ _03266_ _03300_ _03307_ _00284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06231__B _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11985__CLK net438 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09723_ _04436_ _04447_ _04448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06935_ u_cpu.rf_ram_if.rdata1\[0\] u_cpu.rf_ram_if.rtrig1 _02544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_41_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11303__A2 _05547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08937__I _03909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09654_ _04237_ _04384_ _04386_ _00876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_41_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06866_ _01422_ _02466_ _02475_ _02476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_83_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08180__A1 _03415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06885__C _02139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08605_ u_cpu.rf_ram.memory\[143\]\[0\] _03701_ _03702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05817_ u_arbiter.i_wb_cpu_dbus_adr\[4\] _01461_ _01462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09585_ u_arbiter.i_wb_cpu_rdt\[10\] _04334_ _04331_ u_arbiter.i_wb_cpu_dbus_dat\[10\]
+ _04340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06797_ _02401_ _02403_ _02405_ _02407_ _02139_ _02408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_58_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08536_ u_cpu.rf_ram.memory\[73\]\[0\] _03656_ _03657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05748_ _01398_ _01399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06457__I _01803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10814__A1 _05199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08467_ u_cpu.rf_ram.memory\[141\]\[4\] _03613_ _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08483__A2 _03625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11365__CLK net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10290__A2 _04907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07418_ u_cpu.rf_ram.memory\[78\]\[4\] _02929_ _02932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09807__I0 u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08398_ _03570_ u_cpu.rf_ram.memory\[9\]\[4\] _03562_ _03571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07349_ _02881_ _00075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09432__A1 _04140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08235__A2 _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10360_ _02612_ _02640_ u_cpu.cpu.ctrl.i_jump _04954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10042__A2 _02680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09983__A2 _04566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06341__S1 _01841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07994__A1 _03252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09019_ _03957_ _03962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10291_ _04913_ _00986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12030_ _00713_ net312 u_cpu.rf_ram.memory\[91\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06920__I _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09735__A2 _04457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06549__A2 _02162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12863_ u_scanchain_local.clk_out net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12140__CLK net396 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06721__A2 _02332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11058__A1 _05359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11814_ _00510_ net370 u_cpu.rf_ram.memory\[70\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11708__CLK net425 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11745_ _00002_ net252 u_cpu.rf_ram.rdata\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08474__A2 _03610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12290__CLK net501 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11676_ _00380_ net288 u_cpu.rf_ram.memory\[58\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10627_ _05127_ _01108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11858__CLK net420 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09423__A1 u_cpu.rf_ram.memory\[112\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[2\]_CLK net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10033__A2 _04502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11230__A1 _02722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10558_ _05083_ _05088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06332__S1 _01827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout106_I net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10489_ _04813_ _05044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09726__A2 _04450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12228_ _00911_ net360 u_cpu.cpu.immdec.imm30_25\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07737__A1 _03078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12159_ _00842_ net310 u_cpu.rf_ram.memory\[33\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout475_I net476 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06720_ u_cpu.rf_ram.memory\[64\]\[5\] u_cpu.rf_ram.memory\[65\]\[5\] u_cpu.rf_ram.memory\[66\]\[5\]
+ u_cpu.rf_ram.memory\[67\]\[5\] _01798_ _02040_ _02332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_65_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06651_ _02257_ _02259_ _02261_ _02263_ _01835_ _02264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06712__A2 _02323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11049__A1 _05347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11388__CLK net188 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09370_ _04189_ _00789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06582_ _01857_ _02194_ _01859_ _02195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_94_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08321_ u_cpu.rf_ram.memory\[55\]\[7\] _03512_ _03523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08465__A2 _03613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06315__I2 u_cpu.rf_ram.memory\[70\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08252_ u_cpu.rf_ram.memory\[57\]\[1\] _03474_ _03476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10272__A2 _04898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout19_I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07203_ _02777_ _02778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08183_ u_cpu.rf_ram.memory\[60\]\[5\] _03431_ _03435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07134_ _02711_ _02715_ _02716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_14_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10024__A2 _02682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09965__A2 _02703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06779__A2 _02361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07065_ _01430_ _02543_ _02663_ _00008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06016_ _01632_ _01633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_47_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07728__A1 _03060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10262__I _04893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07967_ _02873_ u_cpu.rf_ram.memory\[6\]\[7\] _03288_ _03297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12163__CLK net498 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09706_ _03114_ u_arbiter.i_wb_cpu_rdt\[14\] _04430_ _04431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__11288__A1 u_cpu.rf_ram.memory\[89\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06918_ u_cpu.cpu.state.o_cnt_r\[0\] u_cpu.cpu.state.o_cnt_r\[1\] u_cpu.cpu.state.o_cnt_r\[2\]
+ u_cpu.cpu.state.o_cnt_r\[3\] _02527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_28_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07898_ _03199_ _03242_ _03251_ _00254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09637_ u_arbiter.i_wb_cpu_rdt\[27\] _04293_ _04359_ u_arbiter.i_wb_cpu_dbus_dat\[27\]
+ _04375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_28_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06849_ _01697_ _02458_ _02459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07900__A1 _03227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09568_ _04318_ _04327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08519_ _03593_ _03643_ _03646_ _00480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_70_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09499_ u_cpu.rf_ram.memory\[33\]\[0\] _04271_ _04272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11530_ _00234_ net488 u_cpu.rf_ram.memory\[139\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10263__A2 _04895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08208__A2 _03440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11461_ _00165_ net227 u_cpu.rf_ram.memory\[47\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10412_ _04986_ _01034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11212__A1 _02849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11392_ _00096_ net221 u_cpu.rf_ram.memory\[78\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10343_ _01537_ _04943_ _04938_ u_cpu.cpu.ctrl.o_ibus_adr\[25\] _04944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09708__A2 _04432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10274_ u_cpu.rf_ram.memory\[30\]\[5\] _04898_ _04902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06490__I1 u_cpu.rf_ram.memory\[41\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07719__A1 _01820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12506__CLK net163 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12013_ _00696_ net411 u_cpu.rf_ram.memory\[36\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout480 net483 net480 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_63_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout491 net492 net491 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__06793__I2 u_cpu.rf_ram.memory\[114\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11279__A1 _02899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11530__CLK net488 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08695__A2 _03747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09892__A1 _04255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06250__S0 _01657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xserv_1_568 io_oeb[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__09910__B _04615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08447__A2 _03596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10254__A2 _04888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11728_ _00432_ net136 u_cpu.rf_ram.memory\[9\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06553__S1 _01942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout223_I net229 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11659_ _00363_ net182 u_cpu.rf_ram.memory\[19\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10006__A2 _04548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12036__CLK net284 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11203__A1 _05454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09947__A2 _04629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06630__A1 _02150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06560__I _01788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12186__CLK net497 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08870_ _03826_ _03859_ _03866_ _00611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07186__A2 _02753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07821_ u_cpu.rf_ram.memory\[129\]\[0\] _03205_ _03206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07752_ u_cpu.rf_ram.memory\[17\]\[2\] _03158_ _03159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08135__A1 _03349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06703_ u_cpu.rf_ram.memory\[120\]\[5\] u_cpu.rf_ram.memory\[121\]\[5\] u_cpu.rf_ram.memory\[122\]\[5\]
+ u_cpu.rf_ram.memory\[123\]\[5\] _01674_ _01905_ _02315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_37_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07683_ _02867_ u_cpu.rf_ram.memory\[4\]\[5\] _03101_ _03108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_93_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09883__A1 u_cpu.rf_ram.memory\[114\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09422_ _04154_ _04214_ _04221_ _00809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06697__A1 _02008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06634_ u_cpu.rf_ram.memory\[68\]\[4\] u_cpu.rf_ram.memory\[69\]\[4\] u_cpu.rf_ram.memory\[70\]\[4\]
+ u_cpu.rf_ram.memory\[71\]\[4\] _01779_ _01930_ _02247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_64_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09353_ u_cpu.rf_ram.memory\[121\]\[3\] _04177_ _04179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08438__A2 _03596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06565_ _01564_ _02116_ _02178_ _00003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_33_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08304_ _03512_ _03513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_139_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09284_ _04063_ _04129_ _04134_ _00758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06496_ u_cpu.rf_ram.memory\[36\]\[3\] u_cpu.rf_ram.memory\[37\]\[3\] u_cpu.rf_ram.memory\[38\]\[3\]
+ u_cpu.rf_ram.memory\[39\]\[3\] _01698_ _02109_ _02110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06544__S1 _01930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08235_ u_cpu.rf_ram.memory\[58\]\[2\] _03465_ _03466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08166_ u_cpu.rf_ram.memory\[61\]\[7\] _03406_ _03424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07117_ _02614_ _02703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12529__CLK net276 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10193__S _04849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08097_ u_cpu.rf_ram.memory\[29\]\[7\] _03368_ _03379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08610__A2 _03704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07048_ _02648_ u_cpu.rf_ram.rdata\[2\] _02652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06470__I _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09781__I _04502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11553__CLK net241 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08374__A1 _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08999_ _03945_ _03950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06924__A2 u_cpu.cpu.bufreg.i_sh_signed vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05727__A3 _01377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08397__I _02863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08126__A1 _03340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10961_ _05268_ _05336_ _05338_ _01231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12700_ u_cpu.rf_ram_if.wdata1_r\[4\] net141 u_cpu.rf_ram_if.wdata1_r\[3\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10892_ u_cpu.rf_ram.memory\[69\]\[5\] _05293_ _05297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12631_ _01310_ net59 u_cpu.rf_ram.memory\[25\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12562_ _01241_ net159 u_cpu.rf_ram.memory\[110\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11513_ _00217_ net320 u_cpu.rf_ram.memory\[119\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12493_ _01172_ net38 u_cpu.rf_ram.memory\[106\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07677__S _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06860__A1 _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09929__A2 _04627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11444_ _00148_ net326 u_cpu.rf_ram.memory\[43\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11375_ _00079_ net122 u_cpu.rf_ram.memory\[7\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06612__A1 _02218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10326_ u_cpu.cpu.ctrl.o_ibus_adr\[17\] _04929_ _04931_ u_cpu.cpu.ctrl.o_ibus_adr\[18\]
+ _04934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_113_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10257_ _04886_ _04890_ _04891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09691__I _04415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09562__B1 _04322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10188_ _04851_ _00945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10172__A1 _04821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06471__S0 _02084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05724__I _01374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08117__A1 _03351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09865__A1 _04497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06223__S0 _01574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06679__A1 _02098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout340_I net345 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09617__A1 u_arbiter.i_wb_cpu_rdt\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout438_I net440 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06350_ _01615_ _01965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_61_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06555__I _01813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09093__A2 _04007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06281_ _01725_ _01896_ _01897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11426__CLK net326 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08840__A2 _03848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08020_ u_cpu.rf_ram.memory\[66\]\[3\] _03328_ _03330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08770__I _03801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11576__CLK net340 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09971_ u_cpu.cpu.immdec.imm30_25\[1\] _04516_ _04667_ _04670_ _04671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_118_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08922_ _03894_ _03896_ _03898_ _00631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_48_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout86_I net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08356__A1 _03501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08211__S _03451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08853_ u_cpu.rf_ram.memory\[131\]\[6\] _03851_ _03856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07804_ _03077_ _03193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_57_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08784_ u_cpu.rf_ram.memory\[134\]\[6\] _03806_ _03811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05996_ _01612_ _01613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08108__A1 u_cpu.rf_ram.memory\[63\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07735_ _03075_ _03142_ _03148_ _00194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06509__I2 u_cpu.rf_ram.memory\[102\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07666_ _03081_ _03091_ _03098_ _00175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08945__I _03915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12201__CLK net384 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09405_ _04200_ u_cpu.rf_ram.memory\[11\]\[7\] _04202_ _04211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_81_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06617_ u_cpu.rf_ram.memory\[112\]\[4\] u_cpu.rf_ram.memory\[113\]\[4\] u_cpu.rf_ram.memory\[114\]\[4\]
+ u_cpu.rf_ram.memory\[115\]\[4\] _02133_ _01908_ _02230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_59_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07597_ _02980_ _03048_ _03050_ _00154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09336_ _04152_ _04161_ _04168_ _00776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06548_ u_cpu.rf_ram.memory\[76\]\[3\] u_cpu.rf_ram.memory\[77\]\[3\] u_cpu.rf_ram.memory\[78\]\[3\]
+ u_cpu.rf_ram.memory\[79\]\[3\] _02047_ _01803_ _02162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_21_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09084__A2 _04004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06517__S1 _01905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07095__A1 _02680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09267_ u_cpu.rf_ram.memory\[34\]\[4\] _04121_ _04124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08831__A2 _03839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06479_ u_cpu.rf_ram.memory\[48\]\[3\] u_cpu.rf_ram.memory\[49\]\[3\] u_cpu.rf_ram.memory\[50\]\[3\]
+ u_cpu.rf_ram.memory\[51\]\[3\] _01657_ _02092_ _02093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_142_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08680__I _03484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08218_ _03455_ _00370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09198_ u_cpu.cpu.ctrl.i_jump _04038_ _04078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08149_ _03070_ _03412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05809__I _01451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08595__A1 u_cpu.rf_ram.memory\[70\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11160_ u_cpu.rf_ram.memory\[26\]\[2\] _05469_ _05470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10111_ _04650_ _04750_ _04792_ _04459_ _04795_ _04796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_11091_ _05419_ _05420_ _05421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08347__A1 _03485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10042_ _02605_ _02680_ _04735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09395__I0 _04190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09847__A1 _04527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11993_ _00012_ net259 u_cpu.rf_ram_if.rdata0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06205__S0 _01820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10944_ _05328_ _01224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11449__CLK net299 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10875_ _04832_ _05286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12614_ _01293_ net51 u_cpu.rf_ram.memory\[27\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09075__A2 _03995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[64\] u_scanchain_local.module_data_in\[63\] net554 u_arbiter.o_wb_cpu_adr\[26\]
+ net23 u_scanchain_local.module_data_in\[64\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
X_12545_ _01224_ net118 u_cpu.rf_ram.memory\[10\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08822__A2 _03836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11599__CLK net244 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12476_ _01155_ net234 u_cpu.rf_ram.memory\[79\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11427_ _00131_ net420 u_cpu.rf_ram.memory\[51\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08586__A1 u_cpu.rf_ram.memory\[70\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11358_ _00062_ net59 u_cpu.rf_ram.memory\[20\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10309_ _04909_ _04924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06692__S0 _02001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11289_ _02915_ _05536_ _05545_ _01352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08338__A1 _03504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout388_I net392 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05850_ _01483_ _01488_ u_arbiter.o_wb_cpu_adr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10696__A2 _05165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12224__CLK net343 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout555_I net556 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09838__A1 _03118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05781_ _01430_ u_cpu.rf_ram_if.wtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_82_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07520_ _02998_ _02985_ _02999_ _00128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10448__A2 _04503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07451_ _02921_ _02940_ _02953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12374__CLK net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06402_ _02014_ _02016_ _02017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05875__A2 _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07382_ u_cpu.rf_ram.memory\[80\]\[3\] _02901_ _02905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09121_ _02569_ _04026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_17_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06333_ _01947_ _01948_ _01949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08813__A2 _03817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09052_ _03912_ _03984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06264_ u_cpu.rf_ram.memory\[44\]\[1\] u_cpu.rf_ram.memory\[45\]\[1\] u_cpu.rf_ram.memory\[46\]\[1\]
+ u_cpu.rf_ram.memory\[47\]\[1\] _01692_ _01879_ _01880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06824__A1 _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08003_ _03264_ _03312_ _03319_ _00291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06195_ _01581_ _01812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_11_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08577__A1 _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10384__A1 _04830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09954_ _04419_ _04514_ _04560_ _04654_ _04655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_28_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06683__S0 _01721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08329__A1 _03491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08905_ _03821_ _03882_ _03887_ _00625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09885_ u_cpu.rf_ram.memory\[114\]\[4\] _04592_ _04595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08836_ _03832_ _03836_ _03845_ _00598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08767_ _03763_ _03791_ _03800_ _00574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05979_ _01595_ _01596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07718_ _01820_ _03136_ _03137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08698_ _03757_ _03747_ _03758_ _00547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07649_ u_cpu.rf_ram.memory\[47\]\[7\] _03063_ _03088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05866__A2 _01453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06195__I _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10660_ _03286_ _04959_ _05150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11741__CLK net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09057__A2 _03973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09319_ _04156_ _04143_ _04157_ _00770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08804__A2 _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10591_ u_cpu.rf_ram.memory\[28\]\[5\] _05104_ _05108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12330_ _01010_ net504 u_cpu.cpu.ctrl.o_ibus_adr\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06923__I u_cpu.cpu.branch_op vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12261_ _00944_ net491 u_arbiter.i_wb_cpu_dbus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06291__A2 _01906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08568__A1 _03676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11212_ _02849_ _02891_ _05500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__07955__S _03289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12192_ _00875_ net498 u_arbiter.i_wb_cpu_dbus_dat\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput7 net7 io_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_68_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11143_ _02767_ _05458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06674__S0 _01812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10127__A1 _02890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11074_ _05354_ _05404_ _05409_ _01273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10025_ _04713_ _04714_ _04719_ _00914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06426__S0 _01787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10678__A2 _05150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08740__A1 u_cpu.rf_ram.memory\[136\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07543__A2 _03008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12397__CLK net200 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11976_ _00016_ net265 u_cpu.rf_ram_if.rdata1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09296__A2 _03970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10927_ u_cpu.rf_ram.memory\[59\]\[2\] _05318_ _05319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10858_ _05273_ _05270_ _05274_ _01192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout136_I net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10789_ _02937_ _05162_ _05231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09843__I1 u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06806__A1 _02150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12528_ _01207_ net276 u_cpu.rf_ram.memory\[84\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout303_I net304 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12459_ _01138_ net37 u_cpu.rf_ram.memory\[104\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout309 net310 net309 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_99_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07782__A2 _03172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06951_ _01371_ _02559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11614__CLK net239 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05902_ u_cpu.cpu.ctrl.o_ibus_adr\[21\] u_cpu.cpu.ctrl.o_ibus_adr\[20\] u_cpu.cpu.ctrl.o_ibus_adr\[19\]
+ _01516_ _01529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_41_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09670_ _03117_ _04395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10669__A2 _05151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06882_ _01703_ _02491_ _02492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10023__C _02682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08731__A1 u_cpu.rf_ram.memory\[136\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07534__A2 _03007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08621_ _03684_ _03701_ _03710_ _00518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05833_ u_cpu.cpu.ctrl.o_ibus_adr\[8\] _01474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_67_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08552_ _03606_ _03656_ _03665_ _00494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05764_ _01413_ _01414_ u_cpu.rf_ram_if.rtrig0 _01378_ _01415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_78_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11764__CLK net508 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout49_I net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07503_ u_cpu.rf_ram.memory\[44\]\[1\] _02985_ _02988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07298__A1 u_cpu.rf_ram.memory\[20\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11094__A2 _02633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08483_ u_cpu.rf_ram.memory\[140\]\[2\] _03625_ _03626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07434_ u_cpu.rf_ram.memory\[42\]\[0\] _02943_ _02944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06896__I1 u_cpu.rf_ram.memory\[65\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10841__A2 _05257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07365_ _02890_ _02891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_109_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07839__I _03215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09104_ u_cpu.rf_ram.memory\[36\]\[0\] _04016_ _04017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06316_ _01627_ _01932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07296_ u_cpu.rf_ram.memory\[20\]\[5\] _02837_ _02841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09035_ _03971_ _03972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07470__A1 _02916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06247_ _01650_ _01863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06273__A2 _01848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06178_ _01627_ _01795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06899__B _01782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07222__A1 u_cpu.rf_ram.memory\[21\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06656__S0 _01813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09937_ _04549_ _04456_ _04502_ _04506_ _04639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_89_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05784__A1 _01432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09868_ _04420_ _04509_ _04443_ _04574_ _04582_ _04583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08722__A1 u_cpu.rf_ram.memory\[49\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08819_ _03834_ _03836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09799_ _04475_ _04442_ _04519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11830_ _00526_ net146 u_cpu.rf_ram.memory\[14\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11761_ _00457_ net481 u_cpu.rf_ram.memory\[141\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10712_ _05140_ _05176_ _05182_ _01138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11692_ _00396_ net331 u_cpu.rf_ram.memory\[56\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10643_ u_cpu.rf_ram.memory\[101\]\[2\] _05138_ _05139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10574_ _01443_ _05096_ _05097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_122_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10596__A1 _05057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12313_ _00993_ net528 u_cpu.cpu.ctrl.o_ibus_adr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10060__A3 _04490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07685__S _03101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12244_ _00927_ net274 u_cpu.rf_ram.memory\[32\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06647__S0 _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[27\] u_arbiter.i_wb_cpu_rdt\[24\] net547 u_arbiter.i_wb_cpu_dbus_dat\[21\]
+ net13 u_arbiter.i_wb_cpu_rdt\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
X_12175_ _00858_ net386 u_arbiter.i_wb_cpu_dbus_dat\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10899__A2 _02831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07764__A2 _02936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08961__A1 _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11126_ _05445_ _05446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_111_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09913__B _04459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11057_ u_cpu.rf_ram.memory\[87\]\[4\] _05396_ _05399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11787__CLK net350 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09405__S _04202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08713__A1 u_cpu.rf_ram.memory\[49\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07516__A2 _02990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10008_ _04643_ _04699_ _04703_ _04555_ _04704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_114_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10520__A1 _05046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06575__I0 u_cpu.rf_ram.memory\[20\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06590__I3 u_cpu.rf_ram.memory\[59\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06327__I0 u_cpu.rf_ram.memory\[136\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout253_I net254 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11959_ _00655_ net465 u_cpu.rf_ram.memory\[125\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10823__A2 _05245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout420_I net423 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout518_I net519 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10036__B1 _04652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07150_ _02723_ _02731_ _02732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12412__CLK net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10587__A1 u_cpu.rf_ram.memory\[28\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09441__A2 _04226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06101_ u_cpu.rf_ram.memory\[108\]\[0\] u_cpu.rf_ram.memory\[109\]\[0\] u_cpu.rf_ram.memory\[110\]\[0\]
+ u_cpu.rf_ram.memory\[111\]\[0\] _01716_ _01717_ _01718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07081_ _02671_ _02672_ _01411_ _02591_ _02673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_06032_ _01648_ _01649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06638__S0 _02047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12562__CLK net159 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout106 net107 net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout117 net119 net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__08952__A1 _03061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07755__A2 _03154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout128 net129 net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_102_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07983_ u_cpu.rf_ram.memory\[68\]\[5\] _03303_ _03307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout139 net148 net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_25_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09722_ _04446_ _04447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_41_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06934_ u_cpu.rf_ram.rdata\[0\] _02542_ _02543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_112_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[12\]_SE net544 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08704__A1 _03761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07507__A2 _02990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09752__I0 u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09653_ u_cpu.rf_ram.memory\[113\]\[0\] _04385_ _04386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06865_ _02468_ _02470_ _02472_ _02474_ _01733_ _02475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_27_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10511__A1 _04091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08604_ _03699_ _03701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05816_ _01452_ _01461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09584_ u_arbiter.i_wb_cpu_dbus_dat\[11\] _04338_ _04339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06810__S0 _01779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06191__A1 _01790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06796_ _01691_ _02406_ _01709_ _02407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08535_ _03654_ _03656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06581__I3 u_cpu.rf_ram.memory\[27\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05747_ _01397_ _01398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08466_ _03598_ _03609_ _03615_ _00458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08953__I _03921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10814__A2 _05245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07417_ _02904_ _02925_ _02931_ _00093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10196__S _04855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06494__A2 _02106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08397_ _02863_ _03570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_17_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09807__I1 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07348_ _02855_ u_cpu.rf_ram.memory\[7\]\[1\] _02879_ _02881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09432__A2 _04226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06877__S0 _01773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07279_ _01658_ _02719_ _02829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA__07994__A2 _03312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09018_ _03900_ _03958_ _03961_ _00664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10290_ _01444_ _04907_ _04910_ u_cpu.cpu.ctrl.o_ibus_adr\[3\] _04913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_105_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09196__A1 u_cpu.cpu.state.genblk1.misalign_trap_sync_r vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[38\]_CLK net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06629__S0 _01922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06422__B _01782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08943__A1 _03913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06141__C _01757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09499__A2 _04271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06801__S0 _02029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11813_ _00509_ net377 u_cpu.rf_ram.memory\[70\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11058__A2 _05392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09120__A1 _03988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11744_ _00001_ net252 u_cpu.rf_ram.rdata\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10805__A2 _05236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12435__CLK net160 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11675_ _00379_ net325 u_cpu.rf_ram.memory\[58\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10018__B1 _04712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09895__S _01440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10626_ u_arbiter.i_wb_cpu_rdt\[29\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[13\]
+ _05123_ _05127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_70_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10557_ _05044_ _05084_ _05087_ _01078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11230__A2 _05243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06868__S0 _01639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12585__CLK net207 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09694__I _04418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07985__A2 _03303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10488_ _05039_ _05041_ _05043_ _01053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_12227_ _00910_ net360 u_cpu.cpu.immdec.imm30_25\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[35\]_SE net549 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08934__A1 u_cpu.rf_ram.memory\[128\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07737__A2 _03142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12158_ _00841_ net309 u_cpu.rf_ram.memory\[33\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11109_ _05433_ _01284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12089_ _00772_ net401 u_cpu.rf_ram.memory\[118\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout370_I net372 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06650_ _02060_ _02262_ _01644_ _02263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_92_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06173__A1 _01786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11049__A2 _05392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06581_ u_cpu.rf_ram.memory\[24\]\[4\] u_cpu.rf_ram.memory\[25\]\[4\] u_cpu.rf_ram.memory\[26\]\[4\]
+ u_cpu.rf_ram.memory\[27\]\[4\] _01622_ _01642_ _02194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__05920__A1 _01524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09111__A1 u_cpu.rf_ram.memory\[36\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08320_ _03507_ _03514_ _03522_ _00405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09662__A2 _04388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06315__I3 u_cpu.rf_ram.memory\[71\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08251_ _03405_ _03473_ _03475_ _00383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_127_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06720__I0 u_cpu.rf_ram.memory\[64\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07389__I _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07202_ _02776_ _02777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08182_ _03417_ _03427_ _03434_ _00355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07133_ _02578_ _02714_ _02715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07425__A1 _02916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06859__S0 _01721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09965__A3 _02677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06779__A3 _02370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07064_ u_cpu.rf_ram_if.rdata0\[1\] _02662_ _02663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05987__A1 _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06015_ _01623_ _01632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08225__I0 _02873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07728__A2 _03142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05739__A1 u_cpu.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10732__A1 _05140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12308__CLK net523 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09553__B _04311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07966_ _03296_ _00277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08948__I _02776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09705_ _04413_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[14\] _04430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_25_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06917_ _01406_ _02477_ _02526_ _00007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_68_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11288__A2 _05534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07897_ u_cpu.rf_ram.memory\[74\]\[7\] _03240_ _03251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09636_ u_arbiter.i_wb_cpu_dbus_dat\[28\] _04319_ _04374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06848_ u_cpu.rf_ram.memory\[52\]\[7\] u_cpu.rf_ram.memory\[53\]\[7\] u_cpu.rf_ram.memory\[54\]\[7\]
+ u_cpu.rf_ram.memory\[55\]\[7\] _01747_ _01748_ _02458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_55_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08884__S _03872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12458__CLK net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07900__A2 _02982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09567_ _04292_ _04326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05911__A1 _01453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06779_ _01760_ _02361_ _02370_ _02389_ _02390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_82_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08518_ u_cpu.rf_ram.memory\[72\]\[1\] _03644_ _03646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09498_ _04269_ _04271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_93_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09653__A2 _04385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11482__CLK net379 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08449_ _03506_ _03604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_12_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07664__A1 _03078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06711__I0 u_cpu.rf_ram.memory\[92\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11460_ _00164_ net227 u_cpu.rf_ram.memory\[47\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10411_ _04190_ u_cpu.rf_ram.memory\[2\]\[2\] _04983_ _04986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11212__A2 _02891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11391_ _00095_ net190 u_cpu.rf_ram.memory\[78\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[58\]_SE net562 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10342_ _04905_ _04943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_3_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10273_ _04824_ _04894_ _04901_ _00980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_79_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07963__S _03288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09019__I _03957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12012_ _00695_ net411 u_cpu.rf_ram.memory\[36\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08858__I _03858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout470 net471 net470 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout481 net483 net481 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_24_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout492 net493 net492 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_111_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09341__A1 u_cpu.rf_ram.memory\[118\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08144__A2 _03408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06378__I _01702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xserv_1_569 io_oeb[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06250__S1 _01660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11825__CLK net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09644__A2 _04322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11727_ _00431_ net127 u_cpu.rf_ram.memory\[9\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07655__A1 _03060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11658_ _00362_ net181 u_cpu.rf_ram.memory\[19\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11975__CLK net263 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10609_ u_arbiter.i_wb_cpu_rdt\[21\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[5\]
+ _05117_ _05118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_fanout216_I net219 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11589_ _00293_ net253 u_cpu.rf_ram.memory\[67\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08907__A1 _03824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10714__A1 _05142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06769__I0 u_cpu.rf_ram.memory\[40\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07820_ _03203_ _03205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11355__CLK net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07672__I _03101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09707__I0 u_arbiter.i_wb_cpu_rdt\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12600__CLK net378 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07751_ _03153_ _03158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09332__A1 _04147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06702_ _02014_ _02313_ _02314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08135__A2 _03395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06288__I _01671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07682_ _03107_ _00182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09421_ u_cpu.rf_ram.memory\[112\]\[5\] _04217_ _04221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06633_ _02039_ _02245_ _02246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07894__A1 _03195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06697__A2 _02308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09352_ _04147_ _04173_ _04178_ _00782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout31_I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06564_ _02166_ _02177_ _02178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09635__A2 _04322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08303_ _02877_ _03425_ _03512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07646__A1 _03084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09283_ u_cpu.rf_ram.memory\[117\]\[2\] _04133_ _04134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10538__I _05071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06495_ _01667_ _02109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08234_ _03460_ _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_14_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08165_ _03086_ _03423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07116_ u_cpu.cpu.immdec.imm11_7\[1\] _02700_ _02701_ u_cpu.cpu.immdec.imm11_7\[0\]
+ _02702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XANTENNA__07949__A2 _02784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08071__A1 _03347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08096_ _03351_ _03370_ _03378_ _00325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_49_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12130__CLK net405 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07047_ _02647_ _02649_ _02651_ _00015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_47_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10705__A1 _05130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08374__A2 _03549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08998_ _03900_ _03946_ _03949_ _00656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10181__A2 _02699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07949_ _02721_ _02784_ _03286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_28_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09323__A1 _03180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08126__A2 _03394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[1\]_CLK net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06198__I _01706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10960_ u_cpu.rf_ram.memory\[85\]\[0\] _05337_ _05338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09619_ u_arbiter.i_wb_cpu_rdt\[21\] _04311_ _04321_ u_arbiter.i_wb_cpu_dbus_dat\[21\]
+ _04327_ u_arbiter.i_wb_cpu_dbus_dat\[22\] _04363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__07885__A1 _03186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06688__A2 _02299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10891_ _05280_ _05289_ _05296_ _01203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_43_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12630_ _01309_ net53 u_cpu.rf_ram.memory\[25\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11998__CLK net400 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12561_ _01240_ net162 u_cpu.rf_ram.memory\[110\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07637__A1 u_cpu.rf_ram.memory\[47\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11512_ _00216_ net319 u_cpu.rf_ram.memory\[119\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12492_ _01171_ net38 u_cpu.rf_ram.memory\[106\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11443_ _00147_ net295 u_cpu.rf_ram.memory\[43\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06860__A2 _02469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08062__A1 _03335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11374_ _00078_ net121 u_cpu.rf_ram.memory\[7\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10325_ _04933_ _01000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10183__I _02602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06612__A2 _02220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11378__CLK net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10256_ u_arbiter.i_wb_cpu_dbus_adr\[2\] _02705_ _04890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09562__A1 u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10187_ u_arbiter.i_wb_cpu_dbus_adr\[4\] u_arbiter.i_wb_cpu_dbus_adr\[3\] _04849_
+ _04851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10172__A2 _04836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06766__I3 u_cpu.rf_ram.memory\[59\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06471__S1 _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08117__A2 _03383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09921__B _04626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06128__A1 _01740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11121__A1 _04494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07876__A1 _03197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06223__S1 _01838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout166_I net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12003__CLK net415 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09617__A2 _04293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05740__I u_cpu.cpu.csr_imm vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout333_I net334 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06280_ u_cpu.rf_ram.memory\[100\]\[1\] u_cpu.rf_ram.memory\[101\]\[1\] u_cpu.rf_ram.memory\[102\]\[1\]
+ u_cpu.rf_ram.memory\[103\]\[1\] _01621_ _01895_ _01896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_30_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout500_I net502 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12153__CLK net310 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08053__A1 u_cpu.rf_ram.memory\[65\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout8 u_arbiter.i_wb_cpu_ack net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10935__A1 u_cpu.rf_ram.memory\[59\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09970_ _04498_ _04668_ _04669_ _04670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_89_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07800__A1 _03188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06603__A2 _02187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08921_ u_cpu.rf_ram.memory\[128\]\[0\] _03897_ _03898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09553__A1 u_arbiter.i_wb_cpu_dbus_dat\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08356__A2 _03537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08852_ _03828_ _03848_ _03855_ _00604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout79_I net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07803_ _03191_ _03183_ _03192_ _00218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06757__I3 u_cpu.rf_ram.memory\[27\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08783_ _03759_ _03803_ _03810_ _00580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05995_ _01581_ _01612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08108__A2 _03386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07734_ u_cpu.rf_ram.memory\[16\]\[3\] _03146_ _03148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11112__A1 _02566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07665_ u_cpu.rf_ram.memory\[50\]\[5\] _03094_ _03098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09404_ _04210_ _00802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06616_ _01904_ _02228_ _01679_ _02229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_55_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07596_ u_cpu.rf_ram.memory\[48\]\[0\] _03049_ _03050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09335_ u_cpu.rf_ram.memory\[118\]\[4\] _04165_ _04168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06547_ _01797_ _02160_ _02161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07095__A2 _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09266_ _04066_ _04117_ _04123_ _00751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06478_ _01659_ _02092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08217_ _02861_ u_cpu.rf_ram.memory\[5\]\[3\] _03451_ _03455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08419__I0 _03570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09197_ _03111_ _04027_ _04076_ _04077_ _00727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_107_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06481__I _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08148_ _03410_ _03407_ _03411_ _00344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11520__CLK net430 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08595__A2 _03691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08079_ _03367_ _02967_ _03368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10110_ _04397_ _04794_ _04795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11090_ _01386_ u_cpu.cpu.genblk3.csr.mcause3_0\[1\] _05420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09544__A1 u_arbiter.i_wb_cpu_dbus_dat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08347__A2 _03537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11670__CLK net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10041_ _04732_ _04733_ _04734_ _04467_ _00915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06358__A1 _01630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11992_ _00011_ net259 u_cpu.rf_ram_if.rdata0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12026__CLK net490 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09847__A2 _04456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10943_ _04188_ u_cpu.rf_ram.memory\[10\]\[1\] _05326_ _05328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06205__S1 _01821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10874_ _05284_ _05271_ _05285_ _01197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06530__A1 _01761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09032__I _03893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12176__CLK net387 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12613_ _01292_ net51 u_cpu.rf_ram.memory\[27\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12544_ _01223_ net126 u_cpu.rf_ram.memory\[10\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07086__A2 _02674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10090__A1 _04550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[57\] u_scanchain_local.module_data_in\[56\] net562 u_arbiter.o_wb_cpu_adr\[19\]
+ net31 u_scanchain_local.module_data_in\[57\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__06833__A2 _02442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12475_ _01154_ net232 u_cpu.rf_ram.memory\[79\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08035__A1 _03335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11426_ _00130_ net326 u_cpu.rf_ram.memory\[51\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12045__D _00728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08586__A2 _03688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11357_ _00061_ net56 u_cpu.rf_ram.memory\[20\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10308_ _04923_ _00993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_10_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06692__S1 _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11288_ u_cpu.rf_ram.memory\[89\]\[7\] _05534_ _05545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09535__A1 _04285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08338__A2 _03526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10239_ u_arbiter.i_wb_cpu_dbus_adr\[28\] u_arbiter.i_wb_cpu_dbus_adr\[27\] _04848_
+ _04879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10641__I _04816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05735__I u_cpu.cpu.state.genblk1.misalign_trap_sync_r vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout283_I net284 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05780_ _01401_ _01430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_19_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07950__I _03286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07849__A1 _03191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout450_I net452 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout548_I net549 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07450_ _02916_ _02943_ _02952_ _00105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_78_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06521__A1 _01746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06401_ u_cpu.rf_ram.memory\[124\]\[2\] u_cpu.rf_ram.memory\[125\]\[2\] u_cpu.rf_ram.memory\[126\]\[2\]
+ u_cpu.rf_ram.memory\[127\]\[2\] _02015_ _01737_ _02016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_34_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07381_ _02903_ _02904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09120_ _03988_ _04016_ _04025_ _00702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06332_ u_cpu.rf_ram.memory\[128\]\[1\] u_cpu.rf_ram.memory\[129\]\[1\] u_cpu.rf_ram.memory\[130\]\[1\]
+ u_cpu.rf_ram.memory\[131\]\[1\] _01826_ _01827_ _01948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__11543__CLK net256 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12669__CLK net286 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09051_ _03982_ _03972_ _03983_ _00675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06263_ _01659_ _01879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06824__A2 _02434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08002_ u_cpu.rf_ram.memory\[67\]\[4\] _03316_ _03319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06380__S0 _01705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07397__I _02915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06194_ _01759_ _01809_ _01810_ _01811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10908__A1 _05275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06132__S0 _01747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10384__A2 _04962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09953_ _04650_ _04510_ _04652_ _04653_ _04654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_89_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06683__S1 _01879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08329__A2 _03525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08904_ u_cpu.rf_ram.memory\[22\]\[2\] _03886_ _03887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12049__CLK net271 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09884_ _04247_ _04588_ _04594_ _00898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07001__A2 u_cpu.cpu.ctrl.i_iscomp vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08835_ u_cpu.rf_ram.memory\[132\]\[7\] _03834_ _03845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06060__I0 u_cpu.rf_ram.memory\[56\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08766_ u_cpu.rf_ram.memory\[135\]\[7\] _03789_ _03800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05978_ _01567_ _01595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07860__I _03228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07717_ _02718_ _03135_ _03136_ _00188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__12199__CLK net398 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08888__I0 _03570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08697_ u_cpu.rf_ram.memory\[137\]\[4\] _03753_ _03758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07648_ _03086_ _03087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08892__S _03871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06409__C _01757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06902__I3 u_cpu.rf_ram.memory\[79\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07579_ _02987_ _03036_ _03039_ _00147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09318_ u_cpu.rf_ram.memory\[120\]\[6\] _04148_ _04157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10590_ _05051_ _05100_ _05107_ _01091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09249_ u_cpu.rf_ram.memory\[35\]\[5\] _04109_ _04113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06815__A2 _02425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06371__S0 _01686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12260_ _00943_ net391 u_cpu.cpu.alu.cmp_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07100__I _02602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11211_ _05462_ _05490_ _05499_ _01320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09765__A1 _04412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12191_ _00874_ net498 u_arbiter.i_wb_cpu_dbus_dat\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10375__A2 _04965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11142_ _05456_ _05446_ _05457_ _01293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06674__S1 _02092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11073_ u_cpu.rf_ram.memory\[88\]\[2\] _05408_ _05409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10127__A2 _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10024_ u_cpu.cpu.immdec.imm7 _02682_ _04674_ _04718_ _04719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_27_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06426__S1 _02040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[2\] net8 net548 u_arbiter.i_wb_cpu_dbus_sel\[0\] net15
+ u_arbiter.i_wb_cpu_rdt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__08740__A2 _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11975_ _00015_ net263 u_cpu.rf_ram_if.rdata1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06386__I _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11566__CLK net341 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10926_ _05313_ _05318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_60_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10857_ u_cpu.rf_ram.memory\[108\]\[1\] _05271_ _05274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07059__A2 _02658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08256__A1 _03412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10788_ _05217_ _05221_ _05230_ _01166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10063__A1 _04553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12527_ _01206_ net339 u_cpu.rf_ram.memory\[69\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout129_I net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06362__S0 _01863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06335__B _01419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12458_ _01137_ net37 u_cpu.rf_ram.memory\[104\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09756__A1 _04468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11409_ _00113_ net224 u_cpu.rf_ram.memory\[46\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12389_ _01068_ net196 u_cpu.rf_ram.memory\[94\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07231__A2 _02796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06665__S1 _01968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout498_I net499 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09508__A1 u_cpu.rf_ram.memory\[33\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06950_ _02556_ _02557_ _02558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input3_I io_in[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05901_ u_cpu.cpu.ctrl.o_ibus_adr\[22\] _01528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_95_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06881_ u_cpu.rf_ram.memory\[112\]\[7\] u_cpu.rf_ram.memory\[113\]\[7\] u_cpu.rf_ram.memory\[114\]\[7\]
+ u_cpu.rf_ram.memory\[115\]\[7\] _02133_ _01699_ _02491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08620_ u_cpu.rf_ram.memory\[143\]\[7\] _03699_ _03710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05832_ _01455_ _01473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11909__CLK net462 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06593__I1 u_cpu.rf_ram.memory\[41\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08551_ u_cpu.rf_ram.memory\[73\]\[7\] _03654_ _03665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05763_ u_cpu.cpu.decode.op26 u_cpu.cpu.decode.co_ebreak _01414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07502_ _02896_ _02987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_74_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08482_ _03620_ _03625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08495__A1 _03285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07298__A2 _02837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07433_ _02941_ _02943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_91_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08247__A1 _03380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07364_ _02716_ _02829_ _02890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08217__S _03451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout8_I u_arbiter.i_wb_cpu_ack vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09103_ _04014_ _04016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06315_ u_cpu.rf_ram.memory\[68\]\[1\] u_cpu.rf_ram.memory\[69\]\[1\] u_cpu.rf_ram.memory\[70\]\[1\]
+ u_cpu.rf_ram.memory\[71\]\[1\] _01792_ _01930_ _01931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_143_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09995__A1 _03115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10054__B2 _04537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07295_ _02763_ _02833_ _02840_ _00062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09034_ _03033_ _03970_ _03971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06246_ _01422_ _01862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06273__A3 _01861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06177_ u_cpu.rf_ram.memory\[68\]\[0\] u_cpu.rf_ram.memory\[69\]\[0\] u_cpu.rf_ram.memory\[70\]\[0\]
+ u_cpu.rf_ram.memory\[71\]\[0\] _01792_ _01793_ _01794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_30_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06105__S0 _01721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06656__S1 _01841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10281__I _04905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08970__A2 _03921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09936_ u_arbiter.i_wb_cpu_rdt\[23\] u_arbiter.i_wb_cpu_rdt\[7\] _01441_ _04638_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10109__A2 u_arbiter.i_wb_cpu_rdt\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06981__A1 u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[9\]_SE net544 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09867_ _04552_ _04582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07525__A3 _02724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08686__I _03490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08818_ _03834_ _03835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11589__CLK net253 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09798_ _04517_ _04518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08749_ _03789_ _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11760_ _00456_ net479 u_cpu.rf_ram.memory\[141\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08486__A1 _03598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10711_ u_cpu.rf_ram.memory\[104\]\[3\] _05180_ _05182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11691_ _00395_ net329 u_cpu.rf_ram.memory\[56\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06887__I2 u_cpu.rf_ram.memory\[94\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10642_ _05131_ _05138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08238__A1 _03415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09986__A1 _04494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10573_ u_arbiter.i_wb_cpu_ack u_arbiter.o_wb_cpu_adr\[1\] _05096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12312_ _00992_ net528 u_cpu.cpu.ctrl.o_ibus_adr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09738__A1 _02616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12243_ _00926_ net480 u_cpu.cpu.genblk3.csr.timer_irq_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07765__I _03165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12174_ _00857_ net363 u_arbiter.i_wb_cpu_dbus_dat\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06647__S1 _01827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12364__CLK net210 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11125_ _05098_ _03033_ _05445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08961__A2 _03922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06972__A1 _01431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11056_ _05357_ _05392_ _05398_ _01266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_42_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09910__A1 _04567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10007_ _04700_ _04702_ _04619_ _04703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08713__A2 _03767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10520__A2 _05060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06575__I1 u_cpu.rf_ram.memory\[21\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11958_ _00654_ net451 u_cpu.rf_ram.memory\[126\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06488__B1 _02097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10909_ u_cpu.rf_ram.memory\[84\]\[3\] _05306_ _05308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout246_I net247 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11889_ _00585_ net470 u_cpu.rf_ram.memory\[133\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10036__A1 _04436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10036__B2 _04608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09977__A1 _04626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10366__I _04958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout413_I net414 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06100_ _01667_ _01717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10587__A2 _05104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07080_ _01370_ _02672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_8_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06031_ _01397_ _01648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07204__A2 _02732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06638__S1 _01793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout107 net108 net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_141_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout118 net119 net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__08952__A2 _03181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout129 net130 net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_07982_ _03264_ _03299_ _03306_ _00283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10034__C _04474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11731__CLK net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09721_ _04438_ _04445_ _04446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06933_ u_cpu.rf_ram.regzero _02542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_60_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09901__A1 _04601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08704__A2 _03748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09652_ _04383_ _04385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06864_ _01766_ _02473_ _01731_ _02474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_fanout61_I net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10511__A2 _02921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05815_ u_cpu.cpu.ctrl.o_ibus_adr\[4\] _01459_ _01460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08603_ _03699_ _03700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09583_ _04318_ _04338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10050__B _04737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06810__S1 _01780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06795_ u_cpu.rf_ram.memory\[116\]\[6\] u_cpu.rf_ram.memory\[117\]\[6\] u_cpu.rf_ram.memory\[118\]\[6\]
+ u_cpu.rf_ram.memory\[119\]\[6\] _02136_ _01707_ _02406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_97_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08534_ _03654_ _03655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05746_ _01390_ _01392_ _01396_ _01397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__08468__A1 _03600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10275__A1 _04827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08465_ u_cpu.rf_ram.memory\[141\]\[3\] _03613_ _03615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07140__A1 _02716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07416_ u_cpu.rf_ram.memory\[78\]\[3\] _02929_ _02931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12237__CLK net359 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08396_ _03569_ _00434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10027__A1 _04404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09968__A1 _03115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07347_ _02880_ _00074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08640__A1 _02937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07443__A2 _02946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07278_ _02778_ _02819_ _02828_ _00057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06877__S1 _01774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09017_ u_cpu.rf_ram.memory\[124\]\[1\] _03959_ _03961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06229_ _01590_ _01844_ _01845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06629__S1 _02151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08943__A2 _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09919_ _04620_ _04622_ _04624_ _04585_ _04625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_24_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06706__A1 _01703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09305__I _04141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06801__S1 _01742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11812_ _00508_ net376 u_cpu.rf_ram.memory\[70\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08459__A1 _03588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10266__A1 _04814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11743_ _00000_ net256 u_cpu.rf_ram.rdata\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07131__A1 u_cpu.cpu.immdec.imm11_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11674_ _00378_ net325 u_cpu.rf_ram.memory\[58\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09959__A1 _04546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10018__B2 _04395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10625_ _05126_ _01107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11604__CLK net243 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10569__A2 _05083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10556_ u_cpu.rf_ram.memory\[96\]\[1\] _05085_ _05087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06868__S1 _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10487_ u_cpu.rf_ram.memory\[97\]\[0\] _05042_ _05043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11754__CLK net490 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09187__A2 _04064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12226_ _00909_ net362 u_cpu.cpu.immdec.imm30_25\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12157_ _00840_ net309 u_cpu.rf_ram.memory\[33\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08934__A2 _03904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11108_ u_cpu.cpu.genblk3.csr.mstatus_mie u_cpu.cpu.genblk3.csr.mstatus_mpie _05415_
+ _05433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_81_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12088_ _00771_ net438 u_cpu.rf_ram.memory\[120\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout196_I net202 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11039_ u_cpu.rf_ram.memory\[111\]\[5\] _05384_ _05388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08698__A1 _03757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout363_I net365 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07370__A1 _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06580_ _01630_ _02192_ _02193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09647__B1 _04329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10257__A1 _04886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout530_I net534 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09111__A2 _04019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06556__S0 _02169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08250_ u_cpu.rf_ram.memory\[57\]\[0\] _03474_ _03475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08870__A1 _03826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06720__I1 u_cpu.rf_ram.memory\[65\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07201_ _02734_ u_cpu.cpu.o_wdata0 _02775_ _02776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_14_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08181_ u_cpu.rf_ram.memory\[60\]\[4\] _03431_ _03434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07132_ _02712_ _01414_ _02713_ _02714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08622__A1 _03285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07425__A2 _02926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09818__C _04395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06859__S1 _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07063_ _01401_ _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05987__A2 _01600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06014_ _01573_ _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09178__A2 _04064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07189__A1 _02734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08925__A2 _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05739__A2 _01389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07965_ _02870_ u_cpu.rf_ram.memory\[6\]\[6\] _03288_ _03296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09704_ _04421_ _04423_ _04428_ _04429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_99_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06916_ _02516_ _02525_ _02526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07896_ _03197_ _03242_ _03250_ _00253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09635_ _04370_ _04322_ _04373_ _00870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_112_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06847_ _02450_ _02452_ _02454_ _02456_ _01784_ _02457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_3_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06795__S0 _02136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09566_ _04324_ _04325_ _00849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06778_ _01422_ _02379_ _02388_ _02389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_58_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10248__A1 u_cpu.cpu.bufreg.i_sh_signed vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05729_ _01373_ _01379_ _01380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08517_ _03588_ _03643_ _03645_ _00479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07113__A1 _01388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09497_ _04269_ _04270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_54_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10799__A2 _05236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06484__I _01671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08448_ _03602_ _03591_ _03603_ _00452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08861__A1 _03813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07664__A2 _03090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08379_ u_cpu.rf_ram.memory\[52\]\[6\] _03553_ _03558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10410_ _04985_ _01033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08613__A1 _03676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11390_ _00094_ net189 u_cpu.rf_ram.memory\[78\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07416__A2 _02929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10341_ _04942_ _01007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_136_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10971__A2 _05340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10272_ u_cpu.rf_ram.memory\[30\]\[4\] _04898_ _04901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12011_ _00694_ net425 u_cpu.rf_ram.memory\[37\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11220__I0 _02860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06927__A1 u_cpu.cpu.decode.opcode\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05991__C _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06242__I3 u_cpu.rf_ram.memory\[27\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout460 net474 net460 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_93_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout471 net472 net471 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout482 net483 net482 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_48_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout493 net494 net493 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_46_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12402__CLK net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09341__A2 _04160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06538__S0 _01922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12552__CLK net212 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11726_ _00430_ net416 u_cpu.rf_ram.memory\[52\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08852__A1 _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07655__A2 _03090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11657_ _00361_ net181 u_cpu.rf_ram.memory\[19\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10608_ _03116_ _05117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_70_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11588_ _00292_ net252 u_cpu.rf_ram.memory\[67\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout111_I net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10539_ u_cpu.rf_ram.memory\[95\]\[2\] _05076_ _05077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10962__A2 _05337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12209_ _00892_ net373 u_cpu.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08907__A2 _03882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10714__A2 _05176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06769__I1 u_cpu.rf_ram.memory\[41\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06997__C _02603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09580__A2 _04329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout480_I net483 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07750_ _03068_ _03154_ _03157_ _00200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09868__B1 _04443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12082__CLK net436 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[22\]_CLK net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10478__A1 _04567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09332__A2 _04161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06701_ u_cpu.rf_ram.memory\[124\]\[5\] u_cpu.rf_ram.memory\[125\]\[5\] u_cpu.rf_ram.memory\[126\]\[5\]
+ u_cpu.rf_ram.memory\[127\]\[5\] _02015_ _01774_ _02313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07681_ _02864_ u_cpu.rf_ram.memory\[4\]\[4\] _03102_ _03107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_77_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06632_ u_cpu.rf_ram.memory\[64\]\[4\] u_cpu.rf_ram.memory\[65\]\[4\] u_cpu.rf_ram.memory\[66\]\[4\]
+ u_cpu.rf_ram.memory\[67\]\[4\] _01798_ _02040_ _02245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09420_ _04152_ _04213_ _04220_ _00808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07894__A2 _03242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06563_ _02168_ _02171_ _02173_ _02176_ _01835_ _02177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_09351_ u_cpu.rf_ram.memory\[121\]\[2\] _04177_ _04178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_u_scanchain_local.scan_flop\[37\]_CLK net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09096__A1 _03984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06529__S0 _02142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06518__B _01744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08302_ _03510_ _03488_ _03511_ _00398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09282_ _04128_ _04133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_fanout24_I net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06494_ _01988_ _02106_ _02107_ _02108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08843__A1 _03819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08233_ _03410_ _03461_ _03464_ _00376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_18_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10650__A1 _05142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08164_ _03421_ _03408_ _03422_ _00349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08225__S _03450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07115_ u_cpu.cpu.immdec.imm11_7\[3\] _02701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08095_ u_cpu.rf_ram.memory\[29\]\[6\] _03373_ _03378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08071__A2 _03356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07046_ _02650_ u_cpu.rf_ram_if.rdata1\[1\] _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08959__I _03921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07957__I0 _02858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10705__A2 _05176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12425__CLK net363 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08997_ u_cpu.rf_ram.memory\[125\]\[1\] _03947_ _03949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06385__A2 _01964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06700__C _01900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07582__A1 _02989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07948_ _02849_ _03285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_84_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09323__A2 _03286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07879_ _03227_ _02938_ _03240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12575__CLK net203 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09618_ _04361_ _04362_ _00864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07885__A2 _03241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10890_ u_cpu.rf_ram.memory\[69\]\[4\] _05293_ _05296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09549_ _04292_ _04311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09087__A1 _03975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12560_ _01239_ net162 u_cpu.rf_ram.memory\[110\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08834__A1 _03830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07637__A2 _03072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11511_ _00215_ net320 u_cpu.rf_ram.memory\[119\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12491_ _01170_ net38 u_cpu.rf_ram.memory\[106\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11442_ _00146_ net295 u_cpu.rf_ram.memory\[43\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11373_ _00077_ net60 u_cpu.rf_ram.memory\[7\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08062__A2 _03356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10324_ u_cpu.cpu.ctrl.o_ibus_adr\[16\] _04929_ _04931_ u_cpu.cpu.ctrl.o_ibus_adr\[17\]
+ _04933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_3_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06073__A1 _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05820__A1 u_cpu.cpu.genblk1.align.ctrl_misal vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10255_ _02591_ _04888_ _04889_ _00974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09011__A1 _03919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09562__A2 _04312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10186_ _04850_ _00944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07573__A1 _03018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06389__I _01595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout290 net306 net290 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_43_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06128__A2 _01743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07876__A2 _03230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09078__A1 _03986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06687__I0 u_cpu.rf_ram.memory\[32\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11709_ _00413_ net416 u_cpu.rf_ram.memory\[54\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout326_I net328 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12689_ u_cpu.rf_ram_if.wdata0_r\[6\] net234 u_cpu.rf_ram_if.wdata0_r\[5\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07948__I _02849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11188__A2 _05481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06439__I0 u_cpu.rf_ram.memory\[136\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09250__A1 _04070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout9 net14 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10935__A2 _05318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11322__CLK net185 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06603__A3 _02196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08920_ _03895_ _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_143_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09002__A1 u_cpu.rf_ram.memory\[125\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08851_ u_cpu.rf_ram.memory\[131\]\[5\] _03851_ _03855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07564__A1 _02994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12598__CLK net279 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07802_ u_cpu.rf_ram.memory\[119\]\[3\] _03189_ _03192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06299__I _01687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05994_ _01610_ _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08782_ u_cpu.rf_ram.memory\[134\]\[5\] _03806_ _03810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07733_ _03071_ _03142_ _03147_ _00193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[48\]_SE net558 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07867__A2 _03233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07664_ _03078_ _03090_ _03097_ _00174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_77_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09403_ _04198_ u_cpu.rf_ram.memory\[11\]\[6\] _04202_ _04210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10871__A1 _05282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06615_ u_cpu.rf_ram.memory\[120\]\[4\] u_cpu.rf_ram.memory\[121\]\[4\] u_cpu.rf_ram.memory\[122\]\[4\]
+ u_cpu.rf_ram.memory\[123\]\[4\] _01674_ _01905_ _02228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_41_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07595_ _03047_ _03049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_41_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06546_ u_cpu.rf_ram.memory\[72\]\[3\] u_cpu.rf_ram.memory\[73\]\[3\] u_cpu.rf_ram.memory\[74\]\[3\]
+ u_cpu.rf_ram.memory\[75\]\[3\] _01934_ _01799_ _02160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09334_ _04150_ _04161_ _04167_ _00775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08816__A1 _03832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06678__I0 u_cpu.rf_ram.memory\[56\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09265_ u_cpu.rf_ram.memory\[34\]\[3\] _04121_ _04123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06477_ _01649_ _02090_ _02091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07858__I _02922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08216_ _03454_ _00369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09196_ u_cpu.cpu.state.genblk1.misalign_trap_sync_r _04038_ _04077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10284__I _04908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08147_ u_cpu.rf_ram.memory\[61\]\[1\] _03408_ _03411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09241__A1 _04061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08078_ _02789_ _03367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05802__A1 _01434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07029_ _02532_ _02633_ _01382_ _01379_ _02634_ _02635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_106_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11815__CLK net477 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08689__I _03493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10040_ u_cpu.cpu.immdec.imm7 _02530_ _04734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07555__A1 _02980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06358__A2 _01972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06002__I _01596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11991_ _00010_ net257 u_cpu.rf_ram_if.rdata0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07307__A1 _02726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10942_ _05327_ _01223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05841__I _01452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10862__A1 _05275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10873_ u_cpu.rf_ram.memory\[108\]\[6\] _05276_ _05285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12612_ _01291_ net51 u_cpu.rf_ram.memory\[27\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08807__A1 _03826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10395__S _04973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12543_ _01222_ net291 u_cpu.rf_ram.memory\[59\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07086__A3 _02677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09480__A1 _04237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06913__S0 _01826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06294__A1 _01746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11345__CLK net217 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10090__A2 _04700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12474_ _01153_ net182 u_cpu.rf_ram.memory\[79\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11425_ _00129_ net291 u_cpu.rf_ram.memory\[44\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08035__A2 _03337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09232__A1 _04072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11356_ _00060_ net56 u_cpu.rf_ram.memory\[20\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11495__CLK net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10307_ u_cpu.cpu.ctrl.o_ibus_adr\[9\] _04922_ _04917_ _01484_ _04923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_125_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11287_ _02912_ _05536_ _05544_ _01351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10238_ _04878_ _00968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10169_ u_cpu.rf_ram.memory\[31\]\[2\] _04840_ _04841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout276_I net280 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12120__CLK net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout443_I net444 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06521__A2 _02134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06400_ _01685_ _02015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_91_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07380_ _02757_ _02903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06331_ _01610_ _01947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06285__A1 _01891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09050_ u_cpu.rf_ram.memory\[123\]\[4\] _03978_ _03983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06262_ _01876_ _01877_ _01878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12270__CLK net530 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08001_ _03262_ _03312_ _03318_ _00290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08026__A2 _03328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11838__CLK net478 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09223__A1 u_cpu.rf_ram.memory\[92\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06193_ _01404_ _01810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_u_scanchain_local.scan_flop\[0\]_CLK net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10908__A2 _05302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08503__S _03633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07785__A1 _03087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06132__S1 _01748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09952_ u_arbiter.i_wb_cpu_rdt\[24\] u_arbiter.i_wb_cpu_rdt\[8\] _01446_ _04653_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout91_I net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08903_ _03881_ _03886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_106_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09883_ u_cpu.rf_ram.memory\[114\]\[3\] _04592_ _04594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10053__B _04737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07537__A1 _02989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08834_ _03830_ _03836_ _03844_ _00597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08765_ _03761_ _03791_ _03799_ _00573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05977_ _01590_ _01593_ _01594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07716_ u_cpu.rf_ram_if.rcnt\[2\] u_cpu.rf_ram_if.rcnt\[1\] _02717_ _03136_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_54_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08696_ _03500_ _03757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_65_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07647_ _02777_ _03086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11368__CLK net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07578_ u_cpu.rf_ram.memory\[43\]\[1\] _03037_ _03039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12613__CLK net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09317_ _03915_ _04156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_70_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06529_ u_cpu.rf_ram.memory\[92\]\[3\] u_cpu.rf_ram.memory\[93\]\[3\] u_cpu.rf_ram.memory\[94\]\[3\]
+ u_cpu.rf_ram.memory\[95\]\[3\] _02142_ _01915_ _02143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_22_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08265__A2 _03472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09248_ _04068_ _04105_ _04112_ _00744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06371__S1 _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10943__S _05326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09179_ _04063_ _04058_ _04065_ _00721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06028__A1 _01637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11021__A1 u_cpu.rf_ram.memory\[86\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11210_ u_cpu.rf_ram.memory\[24\]\[7\] _05488_ _05499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12190_ _00873_ net498 u_arbiter.i_wb_cpu_dbus_dat\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09765__A2 _04486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08413__S _03579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09736__C _04460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07776__A1 u_cpu.rf_ram.memory\[40\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11141_ u_cpu.rf_ram.memory\[27\]\[4\] _05452_ _05457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09308__I _03906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09517__A2 _04034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11072_ _05403_ _05408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07528__A1 _03002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10023_ _04715_ _04716_ _04717_ _02682_ _04718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_7_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12143__CLK net396 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11974_ _00670_ net453 u_cpu.rf_ram.memory\[124\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10835__A1 u_cpu.rf_ram.memory\[83\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10925_ _05273_ _05314_ _05317_ _01216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_17_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07700__A1 u_arbiter.i_wb_cpu_dbus_dat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06354__I2 u_cpu.rf_ram.memory\[18\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10856_ _04813_ _05273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09453__A1 _04237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08256__A2 _03473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10787_ u_cpu.rf_ram.memory\[105\]\[7\] _05219_ _05230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06616__B _01679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10063__A2 _04609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12526_ _01205_ net339 u_cpu.rf_ram.memory\[69\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06362__S1 _01653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08008__A2 _03311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12457_ _01136_ net45 u_cpu.rf_ram.memory\[104\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06019__A1 _01630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09756__A2 _04469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11408_ _00112_ net224 u_cpu.rf_ram.memory\[46\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12388_ _01067_ net196 u_cpu.rf_ram.memory\[94\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11339_ _00043_ net187 u_cpu.rf_ram.memory\[81\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout393_I net394 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05900_ _01524_ _01526_ _01527_ u_arbiter.o_wb_cpu_adr\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06880_ _01672_ _02489_ _01679_ _02490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_45_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08192__A1 u_cpu.rf_ram.memory\[19\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05831_ _01456_ _01471_ _01472_ u_arbiter.o_wb_cpu_adr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout560_I net563 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11079__A1 u_cpu.rf_ram.memory\[88\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05762_ _01412_ _01377_ _01413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08550_ _03604_ _03656_ _03664_ _00493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_78_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11510__CLK net301 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07501_ _02980_ _02984_ _02986_ _00122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08481_ _03593_ _03621_ _03624_ _00464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08495__A2 _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07432_ _02941_ _02942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08792__I _03815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07363_ _02888_ _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08247__A2 _03020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11660__CLK net188 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06258__A1 _01672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09102_ _04014_ _04015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10054__A2 _04738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06314_ _01632_ _01930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_17_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09995__A2 u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07294_ u_cpu.rf_ram.memory\[20\]\[4\] _02837_ _02840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06245__C _01428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09033_ _03180_ _03970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06245_ _01851_ _01854_ _01856_ _01860_ _01428_ _01861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__09837__B _04553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06176_ _01632_ _01793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06105__S1 _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09128__I u_cpu.cpu.mem_bytecnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09935_ _04635_ _04629_ _04637_ _04586_ _00906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_63_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12166__CLK net391 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09866_ _04426_ _04561_ _04581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08817_ _02830_ _03814_ _03834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09797_ _04415_ _04418_ _04517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08748_ _02876_ _03698_ _03789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09683__A1 _04403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08486__A2 _03621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08679_ _03684_ _03735_ _03744_ _00542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10710_ _05137_ _05176_ _05181_ _01137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11690_ _00394_ net331 u_cpu.rf_ram.memory\[56\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06887__I3 u_cpu.rf_ram.memory\[95\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10641_ _04816_ _05137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08238__A2 _03461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06249__A1 _01649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11242__A1 u_cpu.rf_ram.memory\[98\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10572_ _04713_ _05095_ _01085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09986__A2 _04679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12311_ _00991_ net528 u_cpu.cpu.ctrl.o_ibus_adr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12242_ _00925_ net383 u_cpu.cpu.immdec.imm31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09738__A2 _04396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12509__CLK net170 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12173_ _00856_ net386 u_arbiter.i_wb_cpu_dbus_dat\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11124_ _02739_ _05444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08877__I _02849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11055_ u_cpu.rf_ram.memory\[87\]\[3\] _05396_ _05398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11533__CLK net488 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08174__A1 u_cpu.rf_ram.memory\[60\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12659__CLK net160 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10006_ _04701_ _04548_ _04615_ _04612_ _04702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_37_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06575__I2 u_cpu.rf_ram.memory\[22\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06280__S0 _01621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09702__S _04417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10808__A1 _05217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11957_ _00653_ net441 u_cpu.rf_ram.memory\[126\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11683__CLK net324 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06327__I2 u_cpu.rf_ram.memory\[138\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06488__A1 _02091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10908_ _05275_ _05302_ _05307_ _01209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11888_ _00584_ net456 u_cpu.rf_ram.memory\[133\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout141_I net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09426__A1 _04158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10839_ _05206_ _05257_ _05262_ _01185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout239_I net240 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12039__CLK net285 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10036__A2 _04510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11233__A1 u_cpu.rf_ram.memory\[98\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07988__A1 _03270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12509_ _01188_ net170 u_cpu.rf_ram.memory\[83\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout406_I net407 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06030_ _01422_ _01647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12189__CLK net497 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout108 net109 net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout119 net120 net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_07981_ u_cpu.rf_ram.memory\[68\]\[4\] _03303_ _03306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09720_ _04443_ _04444_ _04445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06932_ u_cpu.cpu.bufreg2.i_cnt_done _02537_ _02538_ _02540_ _02541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_60_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07691__I _01437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09651_ _04383_ _04384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06863_ u_cpu.rf_ram.memory\[32\]\[7\] u_cpu.rf_ram.memory\[33\]\[7\] u_cpu.rf_ram.memory\[34\]\[7\]
+ u_cpu.rf_ram.memory\[35\]\[7\] _01767_ _01768_ _02473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_110_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08602_ _03061_ _03698_ _03699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05814_ _01447_ u_cpu.cpu.ctrl.o_ibus_adr\[3\] _01444_ _01459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09582_ _04336_ _04337_ _00853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout54_I net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06794_ _01703_ _02404_ _02405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08533_ _03272_ _03020_ _03654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06100__I _01667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05745_ _01394_ _01395_ _01388_ _01367_ _01396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_58_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08468__A2 _03609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09665__A1 _04251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10275__A2 _04895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08464_ _03595_ _03609_ _03614_ _00457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07415_ _02900_ _02925_ _02930_ _00092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09417__A1 u_cpu.rf_ram.memory\[112\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08395_ _03568_ u_cpu.rf_ram.memory\[9\]\[3\] _03562_ _03569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_52_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10027__A2 u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09968__A2 u_arbiter.i_wb_cpu_rdt\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07346_ _02846_ u_cpu.rf_ram.memory\[7\]\[0\] _02879_ _02880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_143_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11406__CLK net221 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07277_ u_cpu.rf_ram.memory\[18\]\[7\] _02817_ _02828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08640__A2 _03698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07866__I _03228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09016_ _03894_ _03958_ _03960_ _00663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06228_ u_cpu.rf_ram.memory\[4\]\[1\] u_cpu.rf_ram.memory\[5\]\[1\] u_cpu.rf_ram.memory\[6\]\[1\]
+ u_cpu.rf_ram.memory\[7\]\[1\] _01591_ _01592_ _01844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_105_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07087__B _01456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06159_ _01772_ _01775_ _01776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11556__CLK net249 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09918_ _04444_ _04623_ _04624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09849_ _04475_ _04490_ _04565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06706__A2 _02317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11811_ _00507_ net376 u_cpu.rf_ram.memory\[70\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06010__I _01601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08459__A2 _03609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09656__A1 _04242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06945__I _01408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11742_ _00446_ net145 u_cpu.rf_ram.memory\[15\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10266__A2 _04894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11673_ _00377_ net314 u_cpu.rf_ram.memory\[58\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06166__B _01782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10624_ u_arbiter.i_wb_cpu_rdt\[28\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[12\]
+ _05123_ _05126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06890__A1 _01740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12331__CLK net501 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10555_ _05039_ _05084_ _05086_ _01077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06642__A1 _02235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10486_ _05040_ _05042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_scanchain_local.scan_flop\[32\] u_arbiter.i_wb_cpu_rdt\[29\] net549 u_arbiter.i_wb_cpu_dbus_dat\[26\]
+ net16 u_arbiter.i_wb_cpu_rdt\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
X_12225_ _00908_ net359 u_cpu.cpu.immdec.imm24_20\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07198__A2 _02753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09592__B1 _04344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12481__CLK net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12156_ _00839_ net309 u_cpu.rf_ram.memory\[33\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11107_ _05430_ _05431_ _05432_ _02577_ _01283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_96_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12087_ _00770_ net443 u_cpu.rf_ram.memory\[120\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08400__I _02866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11038_ _05359_ _05380_ _05387_ _01259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08698__A2 _03747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout189_I net191 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06253__S0 _01639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07370__A2 _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout356_I net367 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07122__A2 _01372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06556__S1 _01821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11429__CLK net327 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout523_I net527 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08870__A2 _03859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07200_ _02726_ u_cpu.rf_ram_if.wdata1_r\[7\] _02775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_14_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10009__A2 _04667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08180_ _03415_ _03427_ _03433_ _00354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_18_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07131_ u_cpu.cpu.immdec.imm11_7\[1\] _02712_ _02713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08622__A2 _02921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11579__CLK net350 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07062_ _02650_ _02660_ _02661_ _00020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_12_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07681__I0 _02864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06013_ _01398_ _01630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08511__S _03632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06492__S0 _01692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07964_ _03295_ _00276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08138__A1 u_cpu.rf_ram.memory\[62\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09703_ _04425_ _04426_ _04427_ _04428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_96_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06915_ _02518_ _02520_ _02522_ _02524_ _01405_ _02525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_112_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07895_ u_cpu.rf_ram.memory\[74\]\[6\] _03245_ _03250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09886__A1 _04249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09634_ u_arbiter.i_wb_cpu_rdt\[26\] _04290_ _04371_ u_arbiter.i_wb_cpu_dbus_dat\[27\]
+ _04373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_67_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06846_ _01619_ _02455_ _01588_ _02456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_56_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12204__CLK net362 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06795__S1 _01707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09565_ u_arbiter.i_wb_cpu_dbus_dat\[5\] _04295_ _04319_ _03130_ _04325_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06777_ _02381_ _02383_ _02385_ _02387_ _01733_ _02388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_58_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05911__A3 _01535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10248__A2 _02705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08516_ u_cpu.rf_ram.memory\[72\]\[0\] _03644_ _03645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05728_ u_cpu.cpu.decode.opcode\[2\] u_cpu.cpu.branch_op _01379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_09496_ _02803_ _02965_ _04269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07113__A2 _02699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08447_ u_cpu.rf_ram.memory\[142\]\[5\] _03596_ _03603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06172__I0 u_cpu.rf_ram.memory\[64\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08861__A2 _03859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06711__I2 u_cpu.rf_ram.memory\[94\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08378_ _03504_ _03550_ _03557_ _00428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07329_ u_cpu.rf_ram_if.wdata0_r\[5\] u_cpu.rf_ram_if.wdata1_r\[5\] _02736_ _02866_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09810__A1 _04518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08613__A2 _03700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09810__B2 _04525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06624__A1 _01761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10340_ u_cpu.cpu.ctrl.o_ibus_adr\[23\] _04936_ _04938_ _01537_ _04942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10951__S _05325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10271_ _04821_ _04894_ _04900_ _00979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09574__B1 _04331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12010_ _00693_ net425 u_cpu.rf_ram.memory\[37\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06005__I _01621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08421__S _03578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10750__I _04816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout450 net452 net450 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__08129__A1 _03342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout461 net467 net461 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_47_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout472 net473 net472 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_19_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout483 net484 net483 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__09877__A1 _04237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout494 net507 net494 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_115_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10487__A2 _05042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06786__S1 _01693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08301__A1 u_cpu.rf_ram.memory\[56\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06538__S1 _02151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11725_ _00429_ net418 u_cpu.rf_ram.memory\[52\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08852__A2 _03848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11656_ _00360_ net179 u_cpu.rf_ram.memory\[19\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11721__CLK net452 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09919__C _04585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout90 net91 net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_126_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10607_ _05116_ _01099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09801__A1 _04514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11587_ _00291_ net251 u_cpu.rf_ram.memory\[67\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10538_ _05071_ _05076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11871__CLK net511 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout104_I net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10469_ _05006_ _05023_ _05027_ _01050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09565__B1 _04319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12208_ _00891_ net384 u_cpu.cpu.csr_d_sel vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06918__A2 u_cpu.cpu.state.o_cnt_r\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12139_ _00822_ net398 u_cpu.rf_ram.memory\[115\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12227__CLK net360 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout473_I net474 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09868__A1 _04420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09868__B2 _04574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06700_ _02305_ _02307_ _02309_ _02311_ _01900_ _02312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__06226__S0 _01583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07680_ _03106_ _00181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06631_ _02237_ _02239_ _02241_ _02243_ _01925_ _02244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_53_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12377__CLK net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09350_ _04172_ _04177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06562_ _02060_ _02175_ _01419_ _02176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09096__A2 _04004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06529__S1 _01915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08301_ u_cpu.rf_ram.memory\[56\]\[7\] _03486_ _03511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09281_ _04061_ _04129_ _04132_ _00757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06493_ _01417_ _02107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08843__A2 _03847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09896__I _04454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08232_ u_cpu.rf_ram.memory\[58\]\[1\] _03462_ _03464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10650__A2 _05132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout17_I net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08163_ u_cpu.rf_ram.memory\[61\]\[6\] _03413_ _03422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07114_ u_cpu.cpu.immdec.imm11_7\[2\] _02700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08094_ _03349_ _03370_ _03377_ _00324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06701__S1 _01774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07045_ _02646_ _02650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09020__A2 _03962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06465__S0 _01849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08996_ _03894_ _03946_ _03948_ _00655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07582__A2 _03036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06385__A3 _01976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07947_ _03270_ _03275_ _03284_ _00270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07878_ _03199_ _03230_ _03239_ _00246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08531__A1 u_cpu.rf_ram.memory\[72\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09617_ u_arbiter.i_wb_cpu_rdt\[20\] _04293_ _04359_ u_arbiter.i_wb_cpu_dbus_dat\[20\]
+ _04362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_95_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06829_ _01406_ _02390_ _02439_ _00006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09548_ u_arbiter.i_wb_cpu_rdt\[3\] _04310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__10011__S _01447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06495__I _01667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09479_ u_cpu.rf_ram.memory\[116\]\[0\] _04259_ _04260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08834__A2 _03836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11510_ _00214_ net301 u_cpu.rf_ram.memory\[40\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12490_ _01169_ net38 u_cpu.rf_ram.memory\[106\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11441_ _00145_ net325 u_cpu.rf_ram.memory\[41\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11894__CLK net458 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08598__A1 _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09795__B1 _04500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11372_ _00076_ net110 u_cpu.rf_ram.memory\[7\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10323_ _04932_ _00999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07270__A1 _02758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10254_ _01370_ _04888_ _04889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09011__A2 _03947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10185_ u_arbiter.i_wb_cpu_dbus_adr\[3\] u_arbiter.i_wb_cpu_dbus_adr\[2\] _04849_
+ _04850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_79_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09046__I _03906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07573__A2 _03034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout280 net281 net280 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_134_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout291 net294 net291 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08522__A1 _03595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05887__A2 _01512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07089__A1 _02679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08825__A2 _03839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11708_ _00412_ net425 u_cpu.rf_ram.memory\[54\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06687__I1 u_cpu.rf_ram.memory\[33\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12688_ u_cpu.rf_ram_if.wdata0_r\[5\] net234 u_cpu.rf_ram_if.wdata0_r\[4\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11639_ _00343_ net186 u_cpu.rf_ram.memory\[61\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout221_I net223 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout319_I net320 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08589__A1 u_cpu.rf_ram.memory\[70\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06439__I1 u_cpu.rf_ram.memory\[137\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09250__A2 _04106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10148__A1 _04824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09002__A2 _03950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06447__S0 _02061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08850_ _03826_ _03847_ _03854_ _00603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10699__A2 _05163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10943__I0 _04188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08761__A1 _03757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07801_ _03074_ _03191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_29_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08781_ _03757_ _03802_ _03809_ _00579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_6_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05993_ _01609_ _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07732_ u_cpu.rf_ram.memory\[16\]\[2\] _03146_ _03147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08795__I _03490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11767__CLK net479 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08513__A1 _03272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07663_ u_cpu.rf_ram.memory\[50\]\[4\] _03094_ _03097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09402_ _04209_ _00801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06614_ _02014_ _02226_ _02227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09069__A2 _03995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07594_ _03047_ _03048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09333_ u_cpu.rf_ram.memory\[118\]\[3\] _04165_ _04167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06545_ _01929_ _02158_ _01932_ _02159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08816__A2 _03817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09264_ _04063_ _04117_ _04122_ _00750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06476_ u_cpu.rf_ram.memory\[52\]\[3\] u_cpu.rf_ram.memory\[53\]\[3\] u_cpu.rf_ram.memory\[54\]\[3\]
+ u_cpu.rf_ram.memory\[55\]\[3\] _01863_ _01653_ _02090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09559__C _04319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08215_ _02858_ u_cpu.rf_ram.memory\[5\]\[2\] _03451_ _03454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09195_ _02673_ _02677_ _04076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08146_ _03067_ _03410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09241__A2 _04105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07252__A1 _02763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08077_ _03353_ _03357_ _03366_ _00318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07028_ u_cpu.cpu.decode.opcode\[1\] u_cpu.cpu.decode.opcode\[0\] _02536_ _02634_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10139__A1 u_cpu.rf_ram.memory\[32\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06850__I1 u_cpu.rf_ram.memory\[49\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07004__A1 u_arbiter.i_wb_cpu_ibus_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08752__A1 _03745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08979_ _03933_ _03938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11990_ _00009_ net263 u_cpu.rf_ram_if.rdata0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07307__A2 _02578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07315__S _02852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10941_ _04184_ u_cpu.rf_ram.memory\[10\]\[0\] _05326_ _05327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10862__A2 _05270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10872_ _04829_ _05284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12611_ _01290_ net52 u_cpu.rf_ram.memory\[27\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08807__A2 _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12542_ _01221_ net277 u_cpu.rf_ram.memory\[59\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06818__A1 _02409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09480__A2 _04258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06913__S1 _02174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06294__A2 _01909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07491__A1 _02913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12473_ _01152_ net241 u_cpu.rf_ram.memory\[79\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[21\]_CLK net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12072__CLK net284 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11424_ _00128_ net292 u_cpu.rf_ram.memory\[44\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10378__A1 _04821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07243__A1 _02740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11355_ _00059_ net68 u_cpu.rf_ram.memory\[20\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10306_ _04905_ _04922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08991__A1 _03919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11286_ u_cpu.rf_ram.memory\[89\]\[6\] _05539_ _05544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[36\]_CLK net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06621__C _02139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10237_ u_arbiter.i_wb_cpu_dbus_adr\[27\] u_arbiter.i_wb_cpu_dbus_adr\[26\] _04873_
+ _04878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08743__A1 _03759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07546__A2 _03006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10168_ _04835_ _04840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10550__A1 _05057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10099_ _04548_ _04565_ _04550_ _04785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09299__A2 _04143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout171_I net172 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06357__I0 u_cpu.rf_ram.memory\[28\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10302__A1 u_cpu.cpu.ctrl.o_ibus_adr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout269_I net540 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout436_I net442 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06330_ _01819_ _01945_ _01823_ _01946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09471__A2 _04245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06285__A2 _01894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06261_ u_cpu.rf_ram.memory\[40\]\[1\] u_cpu.rf_ram.memory\[41\]\[1\] u_cpu.rf_ram.memory\[42\]\[1\]
+ u_cpu.rf_ram.memory\[43\]\[1\] _01686_ _01688_ _01877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_106_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08000_ u_cpu.rf_ram.memory\[67\]\[3\] _03316_ _03318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[20\]_D u_arbiter.i_wb_cpu_rdt\[17\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06192_ _01760_ _01785_ _01808_ _01809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_102_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09223__A2 _04097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07234__A1 _02773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12565__CLK net162 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09951_ _04443_ _04652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08902_ _03819_ _03882_ _03885_ _00624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09882_ _04244_ _04588_ _04593_ _00897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout84_I net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[15\]_SE net542 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08734__A1 _03750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07537__A2 _03007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06103__I _01595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08833_ u_cpu.rf_ram.memory\[132\]\[6\] _03839_ _03844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08764_ u_cpu.rf_ram.memory\[135\]\[6\] _03794_ _03799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05976_ u_cpu.rf_ram.memory\[4\]\[0\] u_cpu.rf_ram.memory\[5\]\[0\] u_cpu.rf_ram.memory\[6\]\[0\]
+ u_cpu.rf_ram.memory\[7\]\[0\] _01591_ _01592_ _01593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__05942__I u_cpu.cpu.ctrl.o_ibus_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07715_ _02717_ _03135_ _00187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08695_ _03755_ _03747_ _03756_ _00546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07646_ _03084_ _03065_ _03085_ _00168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10844__A2 _05261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07577_ _02980_ _03036_ _03038_ _00146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_90_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09316_ _04154_ _04143_ _04155_ _00769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06528_ _01685_ _02142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__12095__CLK net408 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09462__A2 _04245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[22\]_SI u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09247_ u_cpu.rf_ram.memory\[35\]\[4\] _04109_ _04112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06459_ _01958_ _02072_ _02073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06520__I0 u_cpu.rf_ram.memory\[112\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[11\]_D u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09178_ u_cpu.rf_ram.memory\[90\]\[2\] _04064_ _04065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08129_ _03342_ _03394_ _03399_ _00337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06028__A2 _01643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07225__A1 u_cpu.rf_ram.memory\[21\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11021__A2 _05372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09765__A3 _04487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07776__A2 _03172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11140_ _02762_ _05456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_123_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06823__I1 u_cpu.rf_ram.memory\[129\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11932__CLK net333 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10780__A1 _05209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11071_ _05352_ _05404_ _05407_ _01272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08725__A1 _03761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07528__A2 _03005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10022_ _02625_ _04716_ _04717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06948__I _01371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09324__I _04160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11973_ _00669_ net446 u_cpu.rf_ram.memory\[124\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09150__A1 u_cpu.rf_ram.memory\[91\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10924_ u_cpu.rf_ram.memory\[59\]\[1\] _05315_ _05317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12438__CLK net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06354__I3 u_cpu.rf_ram.memory\[19\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10855_ _05268_ _05270_ _05272_ _01191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10786_ _05215_ _05221_ _05229_ _01165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09453__A2 _04239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12525_ _01204_ net345 u_cpu.rf_ram.memory\[69\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07464__A1 _02907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[62\] u_scanchain_local.module_data_in\[61\] net555 u_arbiter.o_wb_cpu_adr\[24\]
+ net22 u_scanchain_local.module_data_in\[62\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XPHY_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06898__S0 _01779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11260__A2 _05527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11462__CLK net297 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[9\]_D u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12456_ _01135_ net45 u_cpu.rf_ram.memory\[104\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09205__A2 _02586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11407_ _00111_ net218 u_cpu.rf_ram.memory\[46\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06019__A2 _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12387_ _01066_ net195 u_cpu.rf_ram.memory\[94\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_u_scanchain_local.scan_flop\[38\]_SE net552 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08403__I _02869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11338_ _00042_ net187 u_cpu.rf_ram.memory\[81\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05778__A1 _01406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09943__B _04553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11269_ _02915_ _05524_ _05533_ _01344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07519__A2 _02990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08716__A1 u_cpu.rf_ram.memory\[49\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11315__A3 u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout386_I net387 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10523__A1 u_cpu.rf_ram.memory\[94\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08192__A2 _03440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05830_ u_arbiter.i_wb_cpu_dbus_adr\[7\] _01461_ _01472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05761_ _01409_ _01411_ _01412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout553_I net557 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06079__B _01695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07500_ u_cpu.rf_ram.memory\[44\]\[0\] _02985_ _02986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08480_ u_cpu.rf_ram.memory\[140\]\[1\] _03622_ _03624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10826__A2 _05249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07431_ _02938_ _02940_ _02941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11805__CLK net347 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07689__I net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07362_ _02739_ _02888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09444__A2 _04230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09101_ _02830_ _02940_ _04014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06313_ _01777_ _01929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06526__C _02139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07455__A1 _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06889__S0 _01741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07293_ _02758_ _02833_ _02839_ _00061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09032_ _03893_ _03969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06244_ _01857_ _01858_ _01859_ _01860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11955__CLK net440 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07207__A1 u_cpu.raddr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06175_ _01572_ _01792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_11_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07758__A2 _03158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10762__A1 _05213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09934_ u_cpu.cpu.immdec.imm24_20\[3\] _04627_ _04636_ _04637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08707__A1 _03763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09865_ _04497_ _04576_ _04579_ _04580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_63_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10514__A1 u_cpu.rf_ram.memory\[94\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08183__A2 _03431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08816_ _03832_ _03817_ _03833_ _00590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09796_ _03118_ _04516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11335__CLK net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06194__A1 _01759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08747_ _03763_ _03779_ _03788_ _00566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05959_ _01575_ _01576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_45_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05941__A1 _01489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08678_ u_cpu.rf_ram.memory\[39\]\[7\] _03733_ _03744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09683__A2 _04407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07694__A1 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06497__A2 _02110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07629_ u_cpu.rf_ram.memory\[47\]\[2\] _03072_ _03073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11485__CLK net376 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10640_ _05135_ _05132_ _05136_ _01112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06436__C _02050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06249__A2 _01864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07446__A1 _02910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10571_ u_cpu.cpu.bufreg.i_sh_signed _04467_ _05095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11242__A2 _05515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09986__A3 _04681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12310_ _00990_ net524 u_cpu.cpu.ctrl.o_ibus_adr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_6_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06008__I _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12241_ _00924_ net260 u_cpu.cpu.immdec.imm19_12_20\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07749__A2 _03155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12172_ _00855_ net386 u_arbiter.i_wb_cpu_dbus_dat\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10753__A1 _05206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11123_ _03111_ u_cpu.cpu.genblk3.csr.timer_irq_r _04806_ _05443_ _01288_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__12110__CLK net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11054_ _05354_ _05392_ _05397_ _01265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10005_ _04505_ _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08174__A2 _03428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12260__CLK net391 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06575__I3 u_cpu.rf_ram.memory\[23\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06280__S1 _01895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09123__A1 _03111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10808__A2 _05233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11956_ _00652_ net453 u_cpu.rf_ram.memory\[126\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10907_ u_cpu.rf_ram.memory\[84\]\[2\] _05306_ _05307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11887_ _00583_ net456 u_cpu.rf_ram.memory\[133\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10838_ u_cpu.rf_ram.memory\[83\]\[2\] _05261_ _05262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11978__CLK net265 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07302__I _02736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07437__A1 _02897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11233__A2 _05512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09938__B _04423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10769_ _03019_ _05162_ _05219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout134_I net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07988__A2 _03300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12508_ _01187_ net162 u_cpu.rf_ram.memory\[83\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10992__A1 _05357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12439_ _01118_ net85 u_cpu.rf_ram.memory\[101\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout301_I net303 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07980_ _03262_ _03299_ _03305_ _00282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout109 net158 net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_45_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06931_ u_cpu.cpu.bufreg2.i_cnt_done u_cpu.cpu.immdec.imm31 _02539_ _02540_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__12603__CLK net374 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09362__A1 _04158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09650_ _02803_ _04224_ _04383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06862_ _01715_ _02471_ _02472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08601_ _03201_ _03698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05813_ _01456_ _01457_ _01458_ u_arbiter.o_wb_cpu_adr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09581_ u_arbiter.i_wb_cpu_rdt\[9\] _04334_ _04331_ u_arbiter.i_wb_cpu_dbus_dat\[9\]
+ _04337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06793_ u_cpu.rf_ram.memory\[112\]\[6\] u_cpu.rf_ram.memory\[113\]\[6\] u_cpu.rf_ram.memory\[114\]\[6\]
+ u_cpu.rf_ram.memory\[115\]\[6\] _02133_ _01699_ _02404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_23_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09114__A1 _03982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08532_ _03606_ _03644_ _03653_ _00486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05744_ u_cpu.cpu.decode.op21 _01381_ _01395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_58_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08509__S _03632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09665__A2 _04385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout47_I net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08463_ u_cpu.rf_ram.memory\[141\]\[2\] _03613_ _03614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07414_ u_cpu.rf_ram.memory\[78\]\[2\] _02929_ _02930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08394_ _02860_ _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_17_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07212__I _02785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07345_ _02878_ _02879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_108_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07979__A2 _03303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07276_ _02773_ _02819_ _02827_ _00056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09015_ u_cpu.rf_ram.memory\[124\]\[0\] _03959_ _03960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06227_ _01580_ _01842_ _01588_ _01843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__12133__CLK net436 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08043__I _03074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06158_ u_cpu.rf_ram.memory\[80\]\[0\] u_cpu.rf_ram.memory\[81\]\[0\] u_cpu.rf_ram.memory\[82\]\[0\]
+ u_cpu.rf_ram.memory\[83\]\[0\] _01773_ _01774_ _01775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_105_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06089_ _01658_ _01706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12283__CLK net504 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09917_ _04485_ _04601_ _04433_ _04599_ _04520_ _04608_ _04623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XFILLER_28_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09848_ _04545_ _04563_ _04564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07903__A2 _03255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10949__S _05326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09779_ _04496_ _04501_ _00886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09105__A1 _03969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11810_ _00506_ net371 u_cpu.rf_ram.memory\[70\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08419__S _03579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09656__A2 _04384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07323__S _02852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11741_ _00445_ net140 u_cpu.rf_ram.memory\[15\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07667__A1 u_cpu.rf_ram.memory\[50\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11672_ _00376_ net314 u_cpu.rf_ram.memory\[58\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10623_ _05125_ _01106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07419__A1 _02907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06961__I u_cpu.cpu.bufreg2.i_cnt_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10554_ u_cpu.rf_ram.memory\[96\]\[0\] _05085_ _05086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08092__A1 _03347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10974__A1 _05284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08219__I0 _02864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10483__I _04807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10485_ _05040_ _05041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09049__I _03909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12224_ _00907_ net343 u_cpu.cpu.immdec.imm24_20\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12626__CLK net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09592__A1 u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[25\] u_arbiter.i_wb_cpu_rdt\[22\] net543 u_arbiter.i_wb_cpu_dbus_dat\[19\]
+ net10 u_arbiter.i_wb_cpu_rdt\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
X_12155_ _00838_ net309 u_cpu.rf_ram.memory\[33\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06910__B _01628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11106_ _02693_ _05431_ _05432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_1_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12086_ _00769_ net443 u_cpu.rf_ram.memory\[120\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08147__A2 _03408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11037_ u_cpu.rf_ram.memory\[111\]\[4\] _05384_ _05387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11151__A1 _05462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09647__A2 _04322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout251_I net254 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06705__I0 u_cpu.rf_ram.memory\[112\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11939_ _00635_ net464 u_cpu.rf_ram.memory\[128\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout349_I net355 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11206__A2 _05493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout516_I net520 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09804__C1 _04523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07130_ u_cpu.rf_ram_if.genblk1.wtrig0_r _02712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_9_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08083__A1 _03335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07061_ _02646_ u_cpu.rf_ram_if.rdata1\[6\] _02661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06633__A2 _02245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07830__A1 u_cpu.rf_ram.memory\[129\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06012_ _01619_ _01626_ _01628_ _01629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10717__A1 u_cpu.rf_ram.memory\[104\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08630__I0 _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08798__I _03493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07963_ _02867_ u_cpu.rf_ram.memory\[6\]\[5\] _03288_ _03295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_9_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06492__S1 _01879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09335__A1 u_cpu.rf_ram.memory\[118\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09702_ u_arbiter.i_wb_cpu_rdt\[2\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[2\]
+ _04417_ _04427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06914_ _01570_ _02523_ _01644_ _02524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07894_ _03195_ _03242_ _03249_ _00252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11142__A1 _05456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09633_ _04370_ _04371_ _04372_ _00869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06111__I _01595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06845_ u_cpu.rf_ram.memory\[24\]\[7\] u_cpu.rf_ram.memory\[25\]\[7\] u_cpu.rf_ram.memory\[26\]\[7\]
+ u_cpu.rf_ram.memory\[27\]\[7\] _01622_ _01625_ _02455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09564_ u_arbiter.i_wb_cpu_rdt\[5\] _04312_ _04324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06776_ _01993_ _02386_ _01996_ _02387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_82_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08515_ _03642_ _03644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05727_ u_cpu.cpu.decode.op21 _01373_ _01377_ _01378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XANTENNA__07649__A1 u_cpu.rf_ram.memory\[47\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09495_ _04255_ _04259_ _04268_ _00835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08446_ _03503_ _03602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_24_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06711__I3 u_cpu.rf_ram.memory\[95\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08377_ u_cpu.rf_ram.memory\[52\]\[5\] _03553_ _03557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07328_ _02865_ _00070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08074__A1 u_cpu.rf_ram.memory\[64\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12649__CLK net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09810__A2 _04520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07821__A1 u_cpu.rf_ram.memory\[129\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07259_ _02723_ _02790_ _02817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10270_ u_cpu.rf_ram.memory\[30\]\[3\] _04898_ _04900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09574__A1 u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11673__CLK net314 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08377__A2 _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06388__A1 _01715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06730__B _01404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06927__A3 u_cpu.cpu.decode.opcode\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10252__B _02565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout440 net442 net440 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_63_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09326__A1 u_cpu.rf_ram.memory\[118\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08129__A2 _03394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout451 net452 net451 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_43_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout462 net467 net462 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_24_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout473 net474 net473 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_63_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout484 net494 net484 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07117__I _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout495 net499 net495 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_86_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06021__I _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07888__A1 _03188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05902__A4 _01516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12179__CLK net387 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11724_ _00428_ net426 u_cpu.rf_ram.memory\[52\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06312__A1 _01786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07360__I0 _02873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11655_ _00359_ net179 u_cpu.rf_ram.memory\[19\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfanout80 net83 net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_128_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout91 net92 net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_10606_ u_arbiter.i_wb_cpu_rdt\[20\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[4\]
+ _05111_ _05116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11586_ _00290_ net248 u_cpu.rf_ram.memory\[67\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09801__A2 _04423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10537_ _05044_ _05072_ _05075_ _01070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07812__A1 _03197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10468_ _02700_ _05006_ _05026_ _04516_ _05027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_48_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09565__A1 u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08368__A2 _03550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12207_ _00890_ net385 u_cpu.cpu.decode.co_mem_word vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10399_ _04196_ u_cpu.rf_ram.memory\[3\]\[5\] _04972_ _04979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10175__A2 _04840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12138_ _00821_ net403 u_cpu.rf_ram.memory\[115\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout299_I net304 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12069_ _00752_ net282 u_cpu.rf_ram.memory\[34\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09868__A2 _04509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07027__I u_arbiter.i_wb_cpu_dbus_we vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06226__S1 _01841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07879__A1 _03227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout466_I net467 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06630_ _02150_ _02242_ _02153_ _02243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09242__I _04104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10388__I _04972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06561_ u_cpu.rf_ram.memory\[132\]\[3\] u_cpu.rf_ram.memory\[133\]\[3\] u_cpu.rf_ram.memory\[134\]\[3\]
+ u_cpu.rf_ram.memory\[135\]\[3\] _02061_ _02174_ _02175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_80_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08300_ _03509_ _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09280_ u_cpu.rf_ram.memory\[117\]\[1\] _04130_ _04132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11546__CLK net258 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06303__A1 _01766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06492_ u_cpu.rf_ram.memory\[44\]\[3\] u_cpu.rf_ram.memory\[45\]\[3\] u_cpu.rf_ram.memory\[46\]\[3\]
+ u_cpu.rf_ram.memory\[47\]\[3\] _01692_ _01879_ _02106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_33_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08231_ _03405_ _03461_ _03463_ _00375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06815__B _01770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08056__A1 u_cpu.rf_ram.memory\[65\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08162_ _03083_ _03421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10938__A1 _05286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07113_ _01388_ _02699_ u_cpu.cpu.o_wen1 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_88_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11696__CLK net417 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07803__A1 _03191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08093_ u_cpu.rf_ram.memory\[29\]\[5\] _03373_ _03377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07044_ _02648_ u_cpu.rf_ram.rdata\[1\] _02649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06106__I _01417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08359__A2 _03541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10166__A2 _04837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06465__S1 _01965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08995_ u_cpu.rf_ram.memory\[125\]\[0\] _03947_ _03948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07946_ u_cpu.rf_ram.memory\[75\]\[7\] _03273_ _03284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11115__A1 _04952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07877_ u_cpu.rf_ram.memory\[77\]\[7\] _03228_ _03239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12321__CLK net532 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09616_ u_arbiter.i_wb_cpu_dbus_dat\[21\] _04352_ _04361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06828_ _02429_ _02438_ _02439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05976__S0 _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06709__C _02139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09547_ _04309_ _00846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06759_ _02363_ _02365_ _02367_ _02369_ _01784_ _02370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_70_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09478_ _04257_ _04259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_12_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08429_ _03589_ _03590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08047__A1 u_cpu.rf_ram.memory\[65\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11440_ _00144_ net324 u_cpu.rf_ram.memory\[41\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10929__A1 u_cpu.rf_ram.memory\[59\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08598__A2 _03688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09795__B2 _04514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11371_ _00075_ net114 u_cpu.rf_ram.memory\[7\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10322_ u_cpu.cpu.ctrl.o_ibus_adr\[15\] _04929_ _04931_ u_cpu.cpu.ctrl.o_ibus_adr\[16\]
+ _04932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_101_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06016__I _01632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07270__A2 _02818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10253_ _02690_ _03123_ _04887_ _04888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05855__I _01451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07022__A2 u_cpu.cpu.mem_bytecnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10184_ _04848_ _04849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_59_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11419__CLK net291 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11106__A1 _02693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout270 net271 net270 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__06781__A1 _02117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout281 net290 net281 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_93_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout292 net294 net292 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_19_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08522__A2 _03643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10202__S _04855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11569__CLK net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09062__I _03990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07089__A2 _01434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08286__A1 _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10093__B2 _04779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11707_ _00411_ net427 u_cpu.rf_ram.memory\[54\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12687_ u_cpu.rf_ram_if.wdata0_r\[4\] net232 u_cpu.rf_ram_if.wdata0_r\[3\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08038__A1 _03340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08406__I _02872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11638_ _00342_ net179 u_cpu.rf_ram.memory\[62\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07310__I _02851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09786__A1 _04459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08589__A2 _03691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06439__I2 u_cpu.rf_ram.memory\[138\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11569_ _00273_ net110 u_cpu.rf_ram.memory\[6\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09237__I _04104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06447__S1 _01832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12344__CLK net385 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08761__A2 _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07800_ _03188_ _03183_ _03190_ _00217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08780_ u_cpu.rf_ram.memory\[134\]\[4\] _03806_ _03809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05992_ _01397_ _01609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07731_ _03141_ _03146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09710__A1 _04416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08513__A2 _03166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07662_ _03075_ _03090_ _03096_ _00173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_93_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12494__CLK net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09401_ _04196_ u_cpu.rf_ram.memory\[11\]\[5\] _04202_ _04209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_19_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06613_ u_cpu.rf_ram.memory\[124\]\[4\] u_cpu.rf_ram.memory\[125\]\[4\] u_cpu.rf_ram.memory\[126\]\[4\]
+ u_cpu.rf_ram.memory\[127\]\[4\] _02015_ _01737_ _02226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07593_ _02891_ _03005_ _03047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06544_ u_cpu.rf_ram.memory\[68\]\[3\] u_cpu.rf_ram.memory\[69\]\[3\] u_cpu.rf_ram.memory\[70\]\[3\]
+ u_cpu.rf_ram.memory\[71\]\[3\] _01792_ _01930_ _02158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09332_ _04147_ _04161_ _04166_ _00774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08277__A1 _03491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09263_ u_cpu.rf_ram.memory\[34\]\[2\] _04121_ _04122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06475_ _02080_ _02083_ _02086_ _02088_ _01428_ _02089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_72_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08214_ _03453_ _00368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08029__A1 _03270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09194_ _04074_ _04059_ _04075_ _00726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08145_ _03405_ _03407_ _03409_ _00343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10387__A2 _03310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08076_ u_cpu.rf_ram.memory\[64\]\[7\] _03355_ _03366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07252__A2 _02806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07027_ u_arbiter.i_wb_cpu_dbus_we _02633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_66_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06850__I2 u_cpu.rf_ram.memory\[50\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08201__A1 u_cpu.rf_ram.memory\[19\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08752__A2 _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08978_ _03900_ _03934_ _03937_ _00648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07929_ _03273_ _03274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_91_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10940_ _05325_ _05326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_21_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10871_ _05282_ _05271_ _05283_ _01196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06610__S1 _01693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12610_ _01289_ net52 u_cpu.rf_ram.memory\[27\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07315__I0 _02855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10075__A1 _04407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07331__S _02851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12541_ _01220_ net293 u_cpu.rf_ram.memory\[59\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06374__S0 _01692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07491__A2 _02970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12472_ _01151_ net241 u_cpu.rf_ram.memory\[79\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07130__I u_cpu.rf_ram_if.genblk1.wtrig0_r vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09768__A1 _04489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11423_ _00127_ net292 u_cpu.rf_ram.memory\[44\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06126__S0 _01741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10378__A2 _04961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10622__I0 u_arbiter.i_wb_cpu_rdt\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11354_ _00058_ net67 u_cpu.rf_ram.memory\[20\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07243__A2 _02806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10305_ _04921_ _00992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__12367__CLK net210 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08991__A2 _03935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11285_ _02909_ _05536_ _05543_ _01350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10236_ _04877_ _00967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10167_ _04814_ _04836_ _04839_ _00936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10550__A2 _05073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10098_ _04701_ _04750_ _04444_ _04784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_19_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10302__A2 _04915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06349__C _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout164_I net173 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09520__I _04284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10066__A1 _04721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06809__A2 _02419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout331_I net332 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout429_I net433 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06260_ _01683_ _01876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07482__A2 _02973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07040__I _02645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09759__A1 _02680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06191_ _01790_ _01796_ _01801_ _01806_ _01807_ _01808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_11_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10613__I0 u_arbiter.i_wb_cpu_rdt\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09950_ _04650_ _04452_ _04507_ _04420_ _04564_ _04651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__08982__A2 _03938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08901_ u_cpu.rf_ram.memory\[22\]\[1\] _03883_ _03885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09881_ u_cpu.rf_ram.memory\[114\]\[2\] _04592_ _04593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09931__A1 _04573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08734__A2 _03778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08832_ _03828_ _03836_ _03843_ _00596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10541__A2 _05076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05975_ _01576_ _01592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08763_ _03759_ _03791_ _03798_ _00572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_73_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06060__I3 u_cpu.rf_ram.memory\[59\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11884__CLK net468 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07714_ _03119_ _03134_ _03135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08694_ u_cpu.rf_ram.memory\[137\]\[3\] _03753_ _03756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07645_ u_cpu.rf_ram.memory\[47\]\[6\] _03072_ _03085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07576_ u_cpu.rf_ram.memory\[43\]\[0\] _03037_ _03038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09430__I _04225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10057__A1 _04542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09998__A1 _02530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09315_ u_cpu.rf_ram.memory\[120\]\[5\] _04148_ _04155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06527_ _01423_ _02128_ _02140_ _02141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_40_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10576__I _02789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08046__I _03077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09246_ _04066_ _04105_ _04111_ _00743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06458_ u_cpu.rf_ram.memory\[4\]\[3\] u_cpu.rf_ram.memory\[5\]\[3\] u_cpu.rf_ram.memory\[6\]\[3\]
+ u_cpu.rf_ram.memory\[7\]\[3\] _01959_ _02071_ _02072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08670__A1 u_cpu.rf_ram.memory\[39\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09177_ _04057_ _04064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06389_ _01595_ _02004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10604__I0 u_arbiter.i_wb_cpu_rdt\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08128_ u_cpu.rf_ram.memory\[62\]\[2\] _03398_ _03399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07225__A2 _02796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08059_ _03355_ _03356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11309__A1 _02915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10780__A2 _05220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11070_ u_cpu.rf_ram.memory\[88\]\[1\] _05405_ _05407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10021_ _02675_ _02703_ _02680_ _04716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09922__A1 _02679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08725__A2 _03767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11972_ _00668_ net465 u_cpu.rf_ram.memory\[124\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06339__I1 u_cpu.rf_ram.memory\[9\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10923_ _05268_ _05314_ _05316_ _01215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07161__A1 _02733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06595__S0 _01692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10854_ u_cpu.rf_ram.memory\[108\]\[0\] _05271_ _05272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10048__A1 _04715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09989__A1 _01443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10048__B2 _04557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10486__I _05040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11607__CLK net236 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06347__S0 _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10785_ u_cpu.rf_ram.memory\[105\]\[6\] _05224_ _05229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12524_ _01203_ net346 u_cpu.rf_ram.memory\[69\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07464__A2 _02954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06898__S1 _01780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[55\] u_scanchain_local.module_data_in\[54\] net561 u_arbiter.o_wb_cpu_adr\[17\]
+ net29 u_scanchain_local.module_data_in\[55\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
X_12455_ _01134_ net86 u_cpu.rf_ram.memory\[103\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11757__CLK net512 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11406_ _00110_ net221 u_cpu.rf_ram.memory\[46\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09610__B1 _04344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12386_ _01065_ net195 u_cpu.rf_ram.memory\[94\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08964__A2 _03926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11337_ _00041_ net95 u_cpu.rf_ram.memory\[21\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06975__A1 u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05778__A2 _01419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06204__I _01815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11268_ u_cpu.rf_ram.memory\[100\]\[7\] _05522_ _05533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06290__I3 u_cpu.rf_ram.memory\[123\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09913__A1 _04528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10219_ _04868_ _00959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11199_ _05488_ _05493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10523__A2 _05064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout281_I net290 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout379_I net380 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05760_ _01410_ _01411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout546_I net551 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06586__S0 _01812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07430_ _02939_ _02940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_63_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10039__A1 _02674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07361_ _02887_ _00081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06807__C _01757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12532__CLK net275 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06312_ _01786_ _01927_ _01928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09100_ _03988_ _04004_ _04013_ _00694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_17_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08652__A1 u_cpu.rf_ram.memory\[138\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07455__A2 _02954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07292_ u_cpu.rf_ram.memory\[20\]\[3\] _02837_ _02839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06889__S1 _01742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09031_ _03919_ _03959_ _03968_ _00670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06243_ _01587_ _01859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06174_ _01777_ _01791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09601__B1 _04344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12682__CLK net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08955__A2 _03923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06805__I2 u_cpu.rf_ram.memory\[86\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05769__A2 _01367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09933_ _04481_ _04636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06114__I _01662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06018__I0 u_cpu.rf_ram.memory\[28\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09904__A1 _04546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08707__A2 _03748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09864_ _04518_ _04578_ _04579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06718__A1 _02150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08815_ u_cpu.rf_ram.memory\[133\]\[7\] _03815_ _03833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10080__B _04767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09795_ _04435_ _04495_ _04500_ _04514_ _04515_ _00888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_3207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07391__A1 _02910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08746_ u_cpu.rf_ram.memory\[136\]\[7\] _03777_ _03788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[20\]_CLK net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05958_ u_cpu.raddr\[1\] _01575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12062__CLK net285 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05889_ u_cpu.cpu.ctrl.o_ibus_adr\[19\] _01516_ _01519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_26_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08677_ _03682_ _03735_ _03743_ _00541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07628_ _03063_ _03072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07694__A2 _01433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[35\]_CLK net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07559_ u_cpu.rf_ram.memory\[41\]\[2\] _03026_ _03027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06329__S0 _01820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10570_ _05057_ _05085_ _05094_ _01084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08643__A1 u_cpu.rf_ram.memory\[138\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09229_ u_cpu.rf_ram.memory\[92\]\[5\] _04097_ _04101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12240_ _00923_ net342 u_cpu.cpu.immdec.imm19_12_20\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12171_ _00854_ net386 u_arbiter.i_wb_cpu_dbus_dat\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_101_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08946__A2 _03904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10753__A2 _05201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11122_ _02693_ _04038_ _05443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06024__I _01575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11053_ u_cpu.rf_ram.memory\[87\]\[2\] _05396_ _05397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10004_ _04610_ _04700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12405__CLK net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[0\] net3 net552 u_arbiter.o_wb_cpu_cyc net20 u_cpu.cpu.genblk3.csr.i_mtip
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_37_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05932__A2 _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10269__A1 _04817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11955_ _00651_ net440 u_cpu.rf_ram.memory\[126\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06568__S0 _01583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12555__CLK net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10906_ _05301_ _05306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11886_ _00582_ net458 u_cpu.rf_ram.memory\[134\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10837_ _05256_ _05261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_60_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07437__A2 _02942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10768_ _05217_ _05202_ _05218_ _01158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_125_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06496__I0 u_cpu.rf_ram.memory\[36\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12507_ _01186_ net163 u_cpu.rf_ram.memory\[83\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout127_I net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10699_ u_cpu.rf_ram.memory\[103\]\[7\] _05163_ _05174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10992__A2 _05349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12438_ _01117_ net85 u_cpu.rf_ram.memory\[101\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12369_ _01048_ net351 u_cpu.cpu.immdec.imm11_7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout496_I net499 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06930_ u_cpu.cpu.csr_d_sel u_cpu.cpu.decode.opcode\[2\] u_cpu.cpu.branch_op _02539_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_101_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input1_I io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09362__A2 _04174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06861_ u_cpu.rf_ram.memory\[36\]\[7\] u_cpu.rf_ram.memory\[37\]\[7\] u_cpu.rf_ram.memory\[38\]\[7\]
+ u_cpu.rf_ram.memory\[39\]\[7\] _01716_ _02109_ _02471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA_u_scanchain_local.scan_flop\[12\]_SI u_arbiter.i_wb_cpu_dbus_dat\[6\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08600_ _03684_ _03688_ _03697_ _00510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05812_ u_arbiter.i_wb_cpu_dbus_adr\[3\] _01453_ _01458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09580_ u_arbiter.i_wb_cpu_dbus_dat\[10\] _04329_ _04336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06792_ _01672_ _02402_ _01679_ _02403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05923__A2 _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05743_ u_cpu.cpu.genblk3.csr.o_new_irq u_cpu.cpu.state.genblk1.misalign_trap_sync_r
+ _01393_ _01394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_08531_ u_cpu.rf_ram.memory\[72\]\[7\] _03642_ _03653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11216__S _05501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06818__B _01404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08462_ _03608_ _03613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_63_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07413_ _02924_ _02929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08393_ _03567_ _00433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07344_ _02850_ _02877_ _02878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09822__B1 _04503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10432__A1 _04817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07275_ u_cpu.rf_ram.memory\[18\]\[6\] _02822_ _02827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06731__S0 _01831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06226_ u_cpu.rf_ram.memory\[12\]\[1\] u_cpu.rf_ram.memory\[13\]\[1\] u_cpu.rf_ram.memory\[14\]\[1\]
+ u_cpu.rf_ram.memory\[15\]\[1\] _01583_ _01841_ _01842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_30_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09014_ _03957_ _03959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10075__B _04474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06239__I0 u_cpu.rf_ram.memory\[28\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06157_ _01652_ _01774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09050__A1 u_cpu.rf_ram.memory\[123\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06088_ _01704_ _01705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_28_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09916_ _04484_ _04621_ _04622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09353__A2 _04177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09847_ _04527_ _04456_ _04563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11452__CLK net335 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07364__A1 _02716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12578__CLK net172 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11160__A2 _05469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08994__I _03945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09778_ _02675_ _04482_ _04497_ _04500_ _04501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_3037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08729_ _03777_ _03778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07116__A1 u_cpu.cpu.immdec.imm11_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11740_ _00444_ net143 u_cpu.rf_ram.memory\[15\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[28\]_SE net547 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07403__I _02920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10671__A1 _05140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11671_ _00375_ net314 u_cpu.rf_ram.memory\[58\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10622_ u_arbiter.i_wb_cpu_rdt\[27\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[11\]
+ _05123_ _05125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08616__A1 u_cpu.rf_ram.memory\[143\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07419__A2 _02925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10423__A1 _04091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10553_ _05083_ _05085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08092__A2 _03369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06722__S0 _01779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10974__A2 _05337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08234__I _03460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10484_ _02803_ _04959_ _05040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12223_ _00906_ net343 u_cpu.cpu.immdec.imm24_20\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09041__A1 _03975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09592__A2 _04334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12154_ _00837_ net309 u_cpu.rf_ram.memory\[33\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11105_ _04026_ _02572_ _02579_ _05431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_85_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xu_scanchain_local.scan_flop\[18\] u_arbiter.i_wb_cpu_rdt\[15\] net542 u_arbiter.i_wb_cpu_dbus_dat\[12\]
+ net9 u_arbiter.i_wb_cpu_rdt\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
X_12085_ _00768_ net443 u_cpu.rf_ram.memory\[120\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11036_ _05357_ _05380_ _05386_ _01258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05905__A2 _01512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11945__CLK net444 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07107__A1 _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11938_ _00634_ net463 u_cpu.rf_ram.memory\[128\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11869_ _00565_ net516 u_cpu.rf_ram.memory\[136\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06330__A2 _01945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09804__B1 _04503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09804__C2 _04477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout411_I net412 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout509_I net510 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09280__A1 u_cpu.rf_ram.memory\[117\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08083__A2 _03369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06713__S0 _02029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05768__I _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10965__A2 _05340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07060_ _02542_ u_cpu.rf_ram.rdata\[6\] _02660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11325__CLK net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07830__A2 _03208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06011_ _01627_ _01628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11214__I0 _02845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11475__CLK net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06397__A2 _02011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07962_ _03294_ _00275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09701_ u_arbiter.i_wb_cpu_rdt\[4\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[4\]
+ _04417_ _04426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_60_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09335__A2 _04165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06913_ u_cpu.rf_ram.memory\[132\]\[7\] u_cpu.rf_ram.memory\[133\]\[7\] u_cpu.rf_ram.memory\[134\]\[7\]
+ u_cpu.rf_ram.memory\[135\]\[7\] _01826_ _02174_ _02523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_64_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07893_ u_cpu.rf_ram.memory\[74\]\[5\] _03245_ _03249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09632_ u_arbiter.i_wb_cpu_rdt\[25\] _04326_ _04295_ u_arbiter.i_wb_cpu_dbus_dat\[25\]
+ _04372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_110_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06844_ _01590_ _02453_ _02454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10350__B1 _04945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09563_ _04320_ _04323_ _00848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06775_ u_cpu.rf_ram.memory\[32\]\[6\] u_cpu.rf_ram.memory\[33\]\[6\] u_cpu.rf_ram.memory\[34\]\[6\]
+ u_cpu.rf_ram.memory\[35\]\[6\] _01767_ _01994_ _02386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_58_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08514_ _03642_ _03643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05726_ _01375_ _01376_ _01377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_36_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09494_ u_cpu.rf_ram.memory\[116\]\[7\] _04257_ _04268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08846__A1 _03821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10653__A1 _05144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08445_ _03600_ _03590_ _03601_ _00451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_12_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08376_ _03501_ _03549_ _03556_ _00427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10405__A1 _02723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07327_ _02864_ u_cpu.rf_ram.memory\[1\]\[4\] _02852_ _02865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_17_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10584__I _05099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06283__B _01731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07258_ _02778_ _02807_ _02816_ _00049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07821__A2 _03205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06209_ _01613_ _01826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07189_ _02734_ u_cpu.rf_ram_if.wdata0_r\[5\] _02765_ _02766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__09023__A1 _03907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09574__A2 _04312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06632__I0 u_cpu.rf_ram.memory\[64\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout430 net431 net430 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_63_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10252__C _03123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout441 net442 net441 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout452 net455 net452 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_115_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout463 net466 net463 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout474 net475 net474 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_43_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout485 net487 net485 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_24_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout496 net499 net496 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_19_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07888__A2 _03241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09613__I _04294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08229__I _03460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08837__A1 _03002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10644__A1 _05137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11723_ _00427_ net427 u_cpu.rf_ram.memory\[52\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11348__CLK net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11654_ _00358_ net220 u_cpu.rf_ram.memory\[60\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout70 net71 net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_15_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout81 net83 net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_10605_ _05115_ _01098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout92 net108 net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_11585_ _00289_ net248 u_cpu.rf_ram.memory\[67\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10536_ u_cpu.rf_ram.memory\[95\]\[1\] _05073_ _05075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05823__A1 _01456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10467_ _04692_ _05025_ _05026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12206_ _00889_ net383 u_cpu.cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09565__A2 _04295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10398_ _04978_ _01028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06640__C _02050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12137_ _00820_ net403 u_cpu.rf_ram.memory\[115\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07308__I _02849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12068_ _00751_ net282 u_cpu.rf_ram.memory\[34\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout194_I net231 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11019_ u_cpu.rf_ram.memory\[86\]\[5\] _05372_ _05376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07879__A2 _02938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout361_I net362 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12123__CLK net406 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout459_I net460 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06551__A2 _02155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08828__A1 _03824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06560_ _01788_ _02174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06491_ _01876_ _02104_ _02105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07500__A1 u_cpu.rf_ram.memory\[44\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08230_ u_cpu.rf_ram.memory\[58\]\[0\] _03462_ _03463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08161_ _03419_ _03408_ _03420_ _00348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07112_ _02674_ _02699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11060__A1 _05361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08092_ _03347_ _03369_ _03376_ _00323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05814__A1 _01447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07043_ _02542_ _02648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09005__A1 _03910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07567__A1 u_cpu.rf_ram.memory\[41\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06550__C _02050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08994_ _03945_ _03947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07218__I _02791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07945_ _03268_ _03275_ _03283_ _00269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11115__A2 _02576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06790__A2 _02400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07876_ _03197_ _03230_ _03238_ _00245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09615_ _04358_ _04360_ _00863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10874__A1 _05284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10579__I _05099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06827_ _02431_ _02433_ _02435_ _02437_ _01405_ _02438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_84_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05976__S1 _01592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09546_ u_arbiter.i_wb_cpu_rdt\[2\] _04290_ _04308_ _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08049__I _03080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06758_ _01619_ _02368_ _01588_ _02369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_97_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12616__CLK net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09477_ _04257_ _04258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_24_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06689_ _02294_ _02296_ _02298_ _02300_ _01733_ _02301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_19_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08428_ _02920_ _03202_ _03589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09244__A1 _04063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08359_ u_cpu.rf_ram.memory\[53\]\[6\] _03541_ _03546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11640__CLK net188 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10929__A2 _05318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11051__A1 _05352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09795__A2 _04495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11370_ _00074_ net110 u_cpu.rf_ram.memory\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10321_ _04908_ _04931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06741__B _02352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07329__S _02736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10252_ u_cpu.cpu.state.o_cnt_r\[0\] u_cpu.cpu.state.o_cnt_r\[1\] _02565_ _03123_
+ _04887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__11790__CLK net347 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10183_ _02602_ _04848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_78_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06032__I _01648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout260 net261 net260 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout271 net275 net271 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout282 net283 net282 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_43_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout293 net294 net293 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_47_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05871__I _01452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10489__I _04813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10865__A1 _05278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07730__A1 _03068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12296__CLK net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11290__A1 _02789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11706_ _00410_ net428 u_cpu.rf_ram.memory\[54\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06297__B2 _01912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12686_ u_cpu.rf_ram_if.wdata0_r\[3\] net232 u_cpu.rf_ram_if.wdata0_r\[2\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08038__A2 _03337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09235__A1 _02939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11637_ _00341_ net179 u_cpu.rf_ram.memory\[62\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11042__A1 _05363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11568_ _00272_ net114 u_cpu.rf_ram.memory\[6\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10519_ u_cpu.rf_ram.memory\[94\]\[2\] _05064_ _05065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout207_I net208 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11499_ _00203_ net178 u_cpu.rf_ram.memory\[17\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06072__I1 u_cpu.rf_ram.memory\[41\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05991_ _01579_ _01589_ _01594_ _01604_ _01607_ _01608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_78_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06772__A2 _02382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07730_ _03068_ _03142_ _03145_ _00192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05781__I _01430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11513__CLK net320 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09710__A2 _04419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07661_ u_cpu.rf_ram.memory\[50\]\[3\] _03094_ _03096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09400_ _04208_ _00800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06612_ _02218_ _02220_ _02222_ _02224_ _01900_ _02225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_20_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07592_ _03000_ _03037_ _03046_ _00153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_59_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09331_ u_cpu.rf_ram.memory\[118\]\[2\] _04165_ _04166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06543_ _02039_ _02156_ _02157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11224__S _05500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06826__B _01644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06907__S0 _01831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout22_I net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09262_ _04116_ _04121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11281__A1 _02903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06474_ _01857_ _02087_ _01859_ _02088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_33_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06678__I3 u_cpu.rf_ram.memory\[59\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08213_ _02855_ u_cpu.rf_ram.memory\[5\]\[1\] _03451_ _03453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_14_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08029__A2 _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09226__A1 _04066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09193_ u_cpu.rf_ram.memory\[90\]\[7\] _04057_ _04075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10067__C _04526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08144_ u_cpu.rf_ram.memory\[61\]\[0\] _03408_ _03409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08075_ _03351_ _03357_ _03365_ _00317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05956__I _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09529__A2 _04284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07026_ _02591_ _02629_ _02602_ _02632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_136_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12169__CLK net385 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09872__B _04586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10395__I0 _04192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08977_ u_cpu.rf_ram.memory\[126\]\[1\] _03935_ _03937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07928_ _03272_ _03034_ _03273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10847__A1 _05215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07859_ _03227_ _02967_ _03228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07712__A1 _02605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06366__I2 u_cpu.rf_ram.memory\[62\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10870_ u_cpu.rf_ram.memory\[108\]\[5\] _05276_ _05283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09529_ _04292_ _04284_ _04294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_25_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12540_ _01219_ net293 u_cpu.rf_ram.memory\[59\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_101_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06669__I3 u_cpu.rf_ram.memory\[27\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06374__S1 _01879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12471_ _01150_ net46 u_cpu.rf_ram.memory\[99\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11024__A1 _05365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11422_ _00126_ net291 u_cpu.rf_ram.memory\[44\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09768__A2 _04490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06027__I _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07779__A1 _03078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06126__S1 _01742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11353_ _00057_ net98 u_cpu.rf_ram.memory\[18\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10304_ u_cpu.cpu.ctrl.o_ibus_adr\[8\] _04915_ _04917_ u_cpu.cpu.ctrl.o_ibus_adr\[9\]
+ _04921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_10_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11284_ u_cpu.rf_ram.memory\[89\]\[5\] _05539_ _05543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06841__I3 u_cpu.rf_ram.memory\[19\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10235_ u_arbiter.i_wb_cpu_dbus_adr\[26\] u_arbiter.i_wb_cpu_dbus_adr\[25\] _04873_
+ _04877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_49_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11536__CLK net250 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10166_ u_cpu.rf_ram.memory\[31\]\[1\] _04837_ _04839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07951__A1 _03285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10213__S _04861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10097_ u_arbiter.i_wb_cpu_rdt\[18\] u_arbiter.i_wb_cpu_rdt\[2\] _01442_ _04783_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_75_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11686__CLK net299 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout157_I net158 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09456__A1 _04242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08259__A2 _03477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08503__I0 _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06109__I2 u_cpu.rf_ram.memory\[102\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10999_ _02772_ _05363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_43_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06646__B _01823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10066__A2 _04710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11263__A1 _02906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_108_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09208__A1 _02703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09957__B _04657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12669_ _01348_ net286 u_cpu.rf_ram.memory\[89\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout324_I net325 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11015__A1 u_cpu.rf_ram.memory\[86\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09759__A2 _04482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06190_ _01606_ _01807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_102_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10613__I1 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10682__I _05163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08431__A2 _03591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05776__I _01426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06993__A2 _02599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08900_ _03813_ _03882_ _03884_ _00623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09880_ _04587_ _04592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_48_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07991__I _03311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08195__A1 _03410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12461__CLK net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08831_ u_cpu.rf_ram.memory\[132\]\[5\] _03839_ _03843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08762_ u_cpu.rf_ram.memory\[135\]\[5\] _03794_ _03798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05974_ _01573_ _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07713_ _02597_ _01386_ _02674_ _03133_ _03134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__06400__I _01685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10829__A1 _05217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08693_ _03497_ _03755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07644_ _03083_ _03084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_65_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09711__I _04427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07170__A2 u_cpu.rf_ram_if.wdata0_r\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09447__A1 _04158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07575_ _03035_ _03037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09314_ _03912_ _04154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11254__A1 _02888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06526_ _02130_ _02132_ _02135_ _02138_ _02139_ _02140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_34_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09245_ u_cpu.rf_ram.memory\[35\]\[3\] _04109_ _04111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11409__CLK net224 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06457_ _01803_ _02071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06520__I2 u_cpu.rf_ram.memory\[114\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09176_ _03902_ _04063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06388_ _01715_ _02002_ _02003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06808__I0 u_cpu.rf_ram.memory\[64\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08127_ _03393_ _03398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_120_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06291__B _01744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11559__CLK net257 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08058_ _02891_ _02923_ _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11309__A2 _05548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07009_ _02614_ _02616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_81_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08186__A1 _03421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10020_ u_cpu.cpu.immdec.imm19_12_20\[0\] _04715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_49_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09922__A2 _02703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06736__A2 _02347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11971_ _00667_ net445 u_cpu.rf_ram.memory\[124\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09686__A1 _04404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08489__A2 _03625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10922_ u_cpu.rf_ram.memory\[59\]\[0\] _05315_ _05316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06044__S0 _01657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07161__A2 _02740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06595__S1 _01879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10853_ _05269_ _05271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10048__A2 _04738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11245__A1 _05458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09989__A2 u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10784_ _05213_ _05221_ _05228_ _01164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08110__A1 u_cpu.rf_ram.memory\[63\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07141__I _02722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06347__S1 _01599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12523_ _01202_ net346 u_cpu.rf_ram.memory\[69\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12334__CLK net523 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12454_ _01133_ net85 u_cpu.rf_ram.memory\[103\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11405_ _00109_ net221 u_cpu.rf_ram.memory\[46\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09610__A1 u_arbiter.i_wb_cpu_rdt\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[48\] u_scanchain_local.module_data_in\[47\] net558 u_arbiter.o_wb_cpu_adr\[10\]
+ net26 u_scanchain_local.module_data_in\[48\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
X_12385_ _01064_ net195 u_cpu.rf_ram.memory\[94\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09068__I _03990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12484__CLK net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11336_ _00040_ net98 u_cpu.rf_ram.memory\[21\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06814__I3 u_cpu.rf_ram.memory\[79\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06975__A2 _02547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05778__A3 _01423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11267_ _02912_ _05524_ _05532_ _01343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10218_ u_arbiter.i_wb_cpu_dbus_adr\[18\] u_arbiter.i_wb_cpu_dbus_adr\[17\] _04867_
+ _04868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_45_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11198_ _05449_ _05489_ _05492_ _01314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06727__A2 _02338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10149_ _02766_ _04826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout274_I net275 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06586__S1 _02092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout441_I net442 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_56_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout539_I net540 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10039__A2 _02625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11236__A1 _05449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07360_ _02873_ u_cpu.rf_ram.memory\[7\]\[7\] _02878_ _02887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06095__C _01711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06311_ u_cpu.rf_ram.memory\[64\]\[1\] u_cpu.rf_ram.memory\[65\]\[1\] u_cpu.rf_ram.memory\[66\]\[1\]
+ u_cpu.rf_ram.memory\[67\]\[1\] _01787_ _01788_ _01927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_52_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07291_ _02752_ _02833_ _02838_ _00060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08652__A2 _03726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09030_ u_cpu.rf_ram.memory\[124\]\[7\] _03957_ _03968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06242_ u_cpu.rf_ram.memory\[24\]\[1\] u_cpu.rf_ram.memory\[25\]\[1\] u_cpu.rf_ram.memory\[26\]\[1\]
+ u_cpu.rf_ram.memory\[27\]\[1\] _01640_ _01642_ _01858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_50_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11701__CLK net415 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10118__S _01447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06173_ _01786_ _01789_ _01790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09601__A1 u_arbiter.i_wb_cpu_rdt\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10598__I0 u_arbiter.i_wb_cpu_rdt\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06805__I3 u_cpu.rf_ram.memory\[87\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06966__A2 _02565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09932_ u_cpu.cpu.immdec.imm24_20\[2\] _04635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11851__CLK net508 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06018__I1 u_cpu.rf_ram.memory\[29\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09904__A2 _04609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09863_ _04458_ _04577_ _04578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10361__B _04953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08814_ _03509_ _03832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_u_scanchain_local.scan_flop\[9\]_SI u_arbiter.i_wb_cpu_dbus_dat\[3\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06274__S0 _01716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09794_ _02676_ _04395_ _04515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12207__CLK net385 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07391__A2 _02894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06130__I _01650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08745_ _03761_ _03779_ _03787_ _00565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_6_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05957_ _01573_ _01574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_22_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06026__S0 _01640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10278__A2 _04893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08676_ u_cpu.rf_ram.memory\[39\]\[6\] _03738_ _03743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05888_ _01505_ _01516_ _01517_ _01518_ u_arbiter.o_wb_cpu_adr\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_26_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07143__A2 _02724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08340__A1 _03507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06577__S1 _01968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07627_ _03070_ _03071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12357__CLK net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07558_ _03021_ _03026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_41_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06329__S1 _01821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06509_ u_cpu.rf_ram.memory\[100\]\[3\] u_cpu.rf_ram.memory\[101\]\[3\] u_cpu.rf_ram.memory\[102\]\[3\]
+ u_cpu.rf_ram.memory\[103\]\[3\] _02122_ _01895_ _02123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_107_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07489_ _02910_ _02970_ _02977_ _00119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09228_ _04068_ _04093_ _04100_ _00736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11381__CLK net176 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09159_ u_cpu.rf_ram.memory\[91\]\[4\] _04049_ _04052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06406__A1 _01746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12170_ _00853_ net383 u_arbiter.i_wb_cpu_dbus_dat\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11121_ _04494_ _05442_ _01287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07337__S _02734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11052_ _05391_ _05396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_46_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07906__A1 u_cpu.rf_ram.memory\[76\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10003_ _04642_ _04582_ _04699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_7_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07382__A2 _02901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06040__I _01620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09659__A1 _04244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10269__A2 _04894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11954_ _00650_ net440 u_cpu.rf_ram.memory\[126\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06568__S1 _01841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10905_ _05273_ _05302_ _05305_ _01208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11885_ _00581_ net468 u_cpu.rf_ram.memory\[134\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10836_ _05204_ _05257_ _05260_ _01184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10767_ u_cpu.rf_ram.memory\[79\]\[7\] _05200_ _05218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12506_ _01185_ net163 u_cpu.rf_ram.memory\[83\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10441__A2 _04992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10698_ _05146_ _05165_ _05173_ _01133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12437_ _01116_ net85 u_cpu.rf_ram.memory\[101\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06215__I _01788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12368_ _01047_ net210 u_cpu.rf_ram.memory\[93\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06799__I2 u_cpu.rf_ram.memory\[94\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07070__A1 _01430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11319_ u_cpu.rf_ram_if.rcnt\[1\] _02717_ _05563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_99_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12299_ _00981_ net81 u_cpu.rf_ram.memory\[30\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08430__I _03589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout391_I net392 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09898__A1 _04546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout489_I net493 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06256__S0 _01871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06860_ _01610_ _02469_ _02107_ _02470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08570__A1 u_cpu.rf_ram.memory\[71\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07373__A2 _02894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05811_ u_cpu.cpu.ctrl.o_ibus_adr\[3\] _01448_ _01457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_55_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06791_ u_cpu.rf_ram.memory\[120\]\[6\] u_cpu.rf_ram.memory\[121\]\[6\] u_cpu.rf_ram.memory\[122\]\[6\]
+ u_cpu.rf_ram.memory\[123\]\[6\] _01674_ _01676_ _02402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_114_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08530_ _03604_ _03644_ _03652_ _00485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05742_ _01379_ _01384_ _01393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__10401__S _04972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08322__A1 _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08461_ _03593_ _03609_ _03612_ _00456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08873__A2 _03863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11209__A1 _05460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07412_ _02897_ _02925_ _02928_ _00091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_90_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06884__A1 _01691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08392_ _03566_ u_cpu.rf_ram.memory\[9\]\[2\] _03562_ _03567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07343_ _02876_ _02877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_71_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09822__A1 _04497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10432__A2 _04993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07274_ _02768_ _02819_ _02826_ _00055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06731__S1 _01942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09013_ _03957_ _03958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06225_ _01584_ _01841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06239__I1 u_cpu.rf_ram.memory\[29\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06125__I _01675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06156_ _01685_ _01773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09050__A2 _03978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06939__A2 _02547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06087_ _01571_ _01704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_104_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09915_ _04436_ _04566_ _04523_ _04608_ _04472_ _04621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_8_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09889__A1 u_cpu.rf_ram.memory\[114\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09846_ _04425_ _04561_ _04562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09372__S _04186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08561__A1 _03671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09777_ _04499_ _04500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06989_ _02527_ _02592_ _02595_ _02596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_85_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08728_ _03165_ _03698_ _03777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11747__CLK net253 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07116__A2 _02700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06728__C _02050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08659_ _03684_ _03723_ _03732_ _00534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10120__A1 _04467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10671__A2 _05151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11670_ _00374_ net99 u_cpu.rf_ram.memory\[5\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10621_ _05124_ _01105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09813__A1 _04411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08616__A2 _03704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07675__I0 _02855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10552_ _05083_ _05084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10423__A2 _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06463__C _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06722__S1 _01930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10483_ _04807_ _05039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12222_ _00905_ net351 u_cpu.cpu.immdec.imm24_20\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12153_ _00836_ net310 u_cpu.rf_ram.memory\[33\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06486__S0 _01871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11104_ u_cpu.cpu.genblk3.csr.mcause31 _05430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_12084_ _00767_ net437 u_cpu.rf_ram.memory\[120\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11035_ u_cpu.rf_ram.memory\[111\]\[3\] _05384_ _05386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08552__A1 _03606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06789__S1 _01774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07107__A2 _02695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12672__CLK net288 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10111__A1 _04650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11937_ _00633_ net463 u_cpu.rf_ram.memory\[128\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10111__B2 _04459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08855__A2 _03846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06866__A1 _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08626__S _03712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11868_ _00564_ net517 u_cpu.rf_ram.memory\[136\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10819_ _05206_ _05245_ _05250_ _01177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09804__A1 _04436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout237_I net238 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08607__A2 _03701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11799_ _00495_ net368 u_cpu.rf_ram.memory\[71\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09804__B2 _04521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06618__A1 _01746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06713__S1 _01742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07291__A1 _02752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout404_I net407 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06010_ _01601_ _01627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10178__A1 _04830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07961_ _02864_ u_cpu.rf_ram.memory\[6\]\[4\] _03289_ _03294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[34\]_CLK net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09700_ _04405_ _04310_ _04424_ _04425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_96_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06912_ _01611_ _02521_ _02522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_25_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07892_ _03193_ _03241_ _03248_ _00251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08543__A1 u_cpu.rf_ram.memory\[73\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09631_ _04300_ _04285_ _04371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06843_ u_cpu.rf_ram.memory\[28\]\[7\] u_cpu.rf_ram.memory\[29\]\[7\] u_cpu.rf_ram.memory\[30\]\[7\]
+ u_cpu.rf_ram.memory\[31\]\[7\] _02084_ _01577_ _02453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_55_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06829__B _02439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09562_ u_arbiter.i_wb_cpu_rdt\[4\] _04312_ _04322_ u_arbiter.i_wb_cpu_dbus_dat\[4\]
+ _04323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_83_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09205__B _02553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06774_ _01715_ _02384_ _02385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout52_I net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[49\]_CLK net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08513_ _03272_ _03166_ _03642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05725_ u_cpu.cpu.branch_op _01376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_70_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10102__A1 _04469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09493_ _04253_ _04259_ _04267_ _00834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08846__A2 _03847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11026__I _05379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08444_ u_cpu.rf_ram.memory\[142\]\[4\] _03596_ _03601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10653__A2 _05133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08375_ u_cpu.rf_ram.memory\[52\]\[4\] _03553_ _03556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06609__A1 _02008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05959__I _01575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10405__A2 _02850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07326_ _02863_ _02864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07257_ u_cpu.rf_ram.memory\[81\]\[7\] _02805_ _02816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06208_ _01610_ _01825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07188_ _02748_ u_cpu.rf_ram_if.wdata1_r\[5\] _02765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09023__A2 _03958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06139_ _01751_ _01754_ _01755_ _01756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_133_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07585__A2 _03040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06632__I1 u_cpu.rf_ram.memory\[65\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout420 net423 net420 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout431 net433 net431 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout442 net449 net442 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_115_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout453 net455 net453 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_24_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout464 net466 net464 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_101_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout475 net476 net475 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__12695__CLK net260 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout486 net487 net486 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_74_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09829_ _04450_ _04546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout497 net499 net497 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XFILLER_100_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06396__I0 u_cpu.rf_ram.memory\[96\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05899__A2 _01481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10892__A2 _05293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08837__A2 _03814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11722_ _00426_ net450 u_cpu.rf_ram.memory\[52\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10644__A2 _05132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07350__S _02879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11653_ _00357_ net220 u_cpu.rf_ram.memory\[60\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout60 net61 net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout71 net72 net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_122_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10604_ u_arbiter.i_wb_cpu_rdt\[19\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[3\]
+ _05111_ _05115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12075__CLK net318 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout82 net83 net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_11584_ _00288_ net245 u_cpu.rf_ram.memory\[67\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfanout93 net95 net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_141_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10535_ _05039_ _05072_ _05074_ _01069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07273__A1 u_cpu.rf_ram.memory\[18\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09785__B _04457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10466_ _04446_ _05024_ _05025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_139_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[30\] u_arbiter.i_wb_cpu_rdt\[27\] net547 u_arbiter.i_wb_cpu_dbus_dat\[24\]
+ net17 u_arbiter.i_wb_cpu_rdt\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__07025__A1 _02627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12205_ _00888_ net384 u_cpu.cpu.branch_op vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_87_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10397_ _04194_ u_cpu.rf_ram.memory\[3\]\[4\] _04973_ _04978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_48_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07576__A2 _03037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12136_ _00819_ net438 u_cpu.rf_ram.memory\[122\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11912__CLK net458 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10580__A1 u_cpu.rf_ram.memory\[28\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12067_ _00750_ net282 u_cpu.rf_ram.memory\[34\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08525__A1 u_cpu.rf_ram.memory\[72\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11018_ _05359_ _05368_ _05375_ _01251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout187_I net192 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10883__A2 _05290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06551__A3 _02164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout354_I net355 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08828__A2 _03835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06490_ u_cpu.rf_ram.memory\[40\]\[3\] u_cpu.rf_ram.memory\[41\]\[3\] u_cpu.rf_ram.memory\[42\]\[3\]
+ u_cpu.rf_ram.memory\[43\]\[3\] _01686_ _02103_ _02104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__12418__CLK net264 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07500__A2 _02985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout521_I net522 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08160_ u_cpu.rf_ram.memory\[61\]\[5\] _03413_ _03420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09253__A2 _04104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07111_ _02697_ _02698_ _02696_ _00023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11442__CLK net295 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07264__A1 u_cpu.rf_ram.memory\[18\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11060__A2 _05393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08091_ u_cpu.rf_ram.memory\[29\]\[4\] _03373_ _03376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06311__I0 u_cpu.rf_ram.memory\[64\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07042_ _02646_ _02647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09005__A2 _03946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07016__A1 _02605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[18\]_SE net542 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08993_ _03945_ _03946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10571__A1 u_cpu.cpu.bufreg.i_sh_signed vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07944_ u_cpu.rf_ram.memory\[75\]\[6\] _03278_ _03283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06870__S0 _01657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08516__A1 u_cpu.rf_ram.memory\[72\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07875_ u_cpu.rf_ram.memory\[77\]\[6\] _03233_ _03238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09614_ u_arbiter.i_wb_cpu_rdt\[19\] _04347_ _04359_ u_arbiter.i_wb_cpu_dbus_dat\[19\]
+ _04360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_55_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06826_ _02060_ _02436_ _01644_ _02437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09545_ _04304_ _04306_ _04300_ _04307_ _04308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_97_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06757_ u_cpu.rf_ram.memory\[24\]\[6\] u_cpu.rf_ram.memory\[25\]\[6\] u_cpu.rf_ram.memory\[26\]\[6\]
+ u_cpu.rf_ram.memory\[27\]\[6\] _01622_ _01625_ _02368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_77_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12098__CLK net405 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09476_ _02830_ _04224_ _04257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06688_ _01993_ _02299_ _01996_ _02300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09492__A2 _04262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08427_ _03484_ _03588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_106_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08358_ _03504_ _03538_ _03545_ _00420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09244__A2 _04105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07309_ _02804_ _02850_ _02851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__11051__A2 _05392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08289_ u_cpu.rf_ram.memory\[56\]\[4\] _03495_ _03502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10320_ _04930_ _00998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_106_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10251_ _04882_ _04884_ _04886_ _02691_ _00973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_65_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06313__I _01777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10182_ _02699_ _04086_ _04847_ _00943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10562__A1 _05049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06861__S0 _01716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout250 net255 net250 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout261 net262 net261 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_8_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout272 net273 net272 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_120_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout283 net284 net283 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_47_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout294 net298 net294 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_43_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10865__A2 _05270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07144__I u_cpu.rf_ram_if.genblk1.wtrig0_r vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07730__A2 _03142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05741__A1 _01391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11705_ _00409_ net427 u_cpu.rf_ram.memory\[54\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11465__CLK net226 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12685_ u_cpu.rf_ram_if.wdata0_r\[2\] net140 u_cpu.rf_ram_if.wdata0_r\[1\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11290__A2 _02877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11636_ _00340_ net179 u_cpu.rf_ram.memory\[62\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_u_scanchain_local.scan_flop\[32\]_D u_arbiter.i_wb_cpu_rdt\[29\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09235__A2 _03310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11567_ _00271_ net110 u_cpu.rf_ram.memory\[6\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10518_ _05059_ _05064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_13_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11498_ _00202_ net178 u_cpu.rf_ram.memory\[17\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10449_ _04562_ _04700_ _05008_ _05009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_87_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout102_I net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07549__A2 _02936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08746__A1 u_cpu.rf_ram.memory\[136\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12119_ _00802_ net143 u_cpu.rf_ram.memory\[11\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05990_ _01606_ _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_38_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout471_I net472 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09171__A1 u_cpu.rf_ram.memory\[90\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06604__S0 _02001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07660_ _03071_ _03090_ _03095_ _00172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09710__A3 _04434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06611_ _01728_ _02223_ _01663_ _02224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05732__A1 u_cpu.cpu.decode.op21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07591_ u_cpu.rf_ram.memory\[43\]\[7\] _03035_ _03046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11808__CLK net376 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09330_ _04160_ _04165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07989__I _03002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06542_ u_cpu.rf_ram.memory\[64\]\[3\] u_cpu.rf_ram.memory\[65\]\[3\] u_cpu.rf_ram.memory\[66\]\[3\]
+ u_cpu.rf_ram.memory\[67\]\[3\] _01787_ _02040_ _02156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_33_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06907__S1 _01832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09261_ _04061_ _04117_ _04120_ _00749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07485__A1 _02904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06473_ u_cpu.rf_ram.memory\[24\]\[3\] u_cpu.rf_ram.memory\[25\]\[3\] u_cpu.rf_ram.memory\[26\]\[3\]
+ u_cpu.rf_ram.memory\[27\]\[3\] _01640_ _01642_ _02087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__12390__CLK net200 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08212_ _03452_ _00367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout15_I net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09192_ _03918_ _04074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_u_scanchain_local.scan_flop\[23\]_D u_arbiter.i_wb_cpu_rdt\[20\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08143_ _03406_ _03408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07237__A1 _02716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11033__A2 _05384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06842__B _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08985__A1 _03910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08074_ u_cpu.rf_ram.memory\[64\]\[6\] _03360_ _03365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07025_ _02627_ _02630_ _02631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08737__A1 _03752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10544__A1 _05051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06599__I0 u_cpu.rf_ram.memory\[32\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06212__A2 _01828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06843__S0 _02084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11338__CLK net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08976_ _03894_ _03934_ _03936_ _00647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07927_ _02922_ _03272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09162__A1 _03984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07012__I1 u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07858_ _02922_ _03227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06809_ _02039_ _02419_ _02420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06366__I3 u_cpu.rf_ram.memory\[63\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11488__CLK net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07789_ _02877_ _03181_ _03182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07899__I _03059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09528_ _04292_ _04293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09465__A2 _04245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09459_ u_cpu.rf_ram.memory\[115\]\[2\] _04245_ _04246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12470_ _01149_ net46 u_cpu.rf_ram.memory\[99\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_u_scanchain_local.scan_flop\[14\]_D u_arbiter.i_wb_cpu_rdt\[11\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11421_ _00125_ net297 u_cpu.rf_ram.memory\[44\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07228__A1 _02758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11024__A2 _05369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08976__A1 _03894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07779__A2 _03168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11352_ _00056_ net69 u_cpu.rf_ram.memory\[18\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10303_ _04920_ _00991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__12113__CLK net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11283_ _02906_ _05535_ _05542_ _01349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_49_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08728__A1 _03165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10234_ _04876_ _00966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06043__I _01659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10535__A1 _05039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07400__A1 _02578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10165_ _04808_ _04836_ _04838_ _00935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06834__S0 _01640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07951__A2 _03287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10096_ _04772_ _04780_ _04781_ _04782_ _00922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__05962__A1 _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09153__A1 _03975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10838__A2 _05261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07703__A2 _03123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08900__A1 _03813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09456__A2 _04239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10998_ _05361_ _05350_ _05362_ _01244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11263__A2 _05523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11124__I _02739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06218__I _01405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08634__S _03711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12668_ _01347_ net286 u_cpu.rf_ram.memory\[89\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11015__A2 _05372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11619_ _00323_ net103 u_cpu.rf_ram.memory\[29\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout317_I net322 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12599_ _01278_ net278 u_cpu.rf_ram.memory\[88\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08967__A1 _03913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08433__I _03490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06442__A2 _02056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06293__I2 u_cpu.rf_ram.memory\[114\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08719__A1 _03755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10526__A1 _05053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08195__A2 _03439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08830_ _03826_ _03835_ _03842_ _00595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06825__S0 _02061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05792__I _01438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07942__A2 _03278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08761_ _03757_ _03790_ _03797_ _00571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05973_ _01398_ _01590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09144__A1 _03112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07712_ _02605_ _03131_ _03132_ _02684_ _03133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08692_ _03752_ _03747_ _03754_ _00545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10829__A2 _05246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07643_ _02772_ _03083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06837__B _01795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07574_ _03035_ _03036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_41_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11780__CLK net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09447__A2 _04227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07512__I _02906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09313_ _04152_ _04142_ _04153_ _00768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06525_ _01426_ _02139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__10057__A3 _04746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11254__A2 _05523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09998__A3 _04665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09244_ _04063_ _04105_ _04110_ _00742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06456_ _01580_ _02068_ _02069_ _02070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_72_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12136__CLK net438 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09175_ _04061_ _04058_ _04062_ _00720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06387_ u_cpu.rf_ram.memory\[108\]\[2\] u_cpu.rf_ram.memory\[109\]\[2\] u_cpu.rf_ram.memory\[110\]\[2\]
+ u_cpu.rf_ram.memory\[111\]\[2\] _02001_ _01717_ _02002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__05967__I _01575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08958__A1 _03900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08126_ _03340_ _03394_ _03397_ _00336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06808__I1 u_cpu.rf_ram.memory\[65\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10765__A1 _05215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08057_ _03353_ _03338_ _03354_ _00310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07630__A1 _03071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12286__CLK net502 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07008_ _02613_ _02614_ _02615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09375__S _04186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10517__A1 _05044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08186__A2 _03428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09922__A3 _01377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07933__A2 _03275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08959_ _03921_ _03926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09135__A1 _03112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11970_ _00666_ net445 u_cpu.rf_ram.memory\[124\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09686__A2 u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09902__I _04402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07697__A1 u_cpu.cpu.state.genblk1.misalign_trap_sync_r vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10921_ _05313_ _05315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06044__S1 _01660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10852_ _05269_ _05270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09438__A2 _04230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08497__I0 _03560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11245__A2 _05512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10783_ u_cpu.rf_ram.memory\[105\]\[5\] _05224_ _05228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08110__A2 _03386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12522_ _01201_ net346 u_cpu.rf_ram.memory\[69\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12453_ _01132_ net85 u_cpu.rf_ram.memory\[103\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11404_ _00108_ net221 u_cpu.rf_ram.memory\[46\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11503__CLK net295 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12384_ _01063_ net195 u_cpu.rf_ram.memory\[94\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12629__CLK net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09610__A2 _04347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10756__A1 _05209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11335_ _00039_ net98 u_cpu.rf_ram.memory\[21\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07621__A1 _03060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05778__A4 _01428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11266_ u_cpu.rf_ram.memory\[100\]\[6\] _05527_ _05532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08177__A2 _03431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10217_ _02690_ _04867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__11653__CLK net220 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10224__S _04867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08421__I0 _03572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11197_ u_cpu.rf_ram.memory\[24\]\[1\] _05490_ _05492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11181__A1 _05451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10148_ _04824_ _04810_ _04825_ _00931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10079_ _04407_ _04518_ _04749_ _04552_ _04767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__12009__CLK net425 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout267_I net268 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12159__CLK net310 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11236__A2 _05511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06310_ _01917_ _01919_ _01921_ _01924_ _01925_ _01926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_52_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07290_ u_cpu.rf_ram.memory\[20\]\[2\] _02837_ _02838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10995__A1 _05359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06241_ _01596_ _01857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_15_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06172_ u_cpu.rf_ram.memory\[64\]\[0\] u_cpu.rf_ram.memory\[65\]\[0\] u_cpu.rf_ram.memory\[66\]\[0\]
+ u_cpu.rf_ram.memory\[67\]\[0\] _01787_ _01788_ _01789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_8_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09601__A2 _04347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07612__A1 _03000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09931_ _04573_ _04634_ _00905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05736__B _01385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09862_ _04563_ _04568_ _04577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout82_I net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11172__A1 _05098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08813_ _03830_ _03817_ _03831_ _00589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06411__I _01565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06274__S1 _01717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09793_ _04421_ _04514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09117__A1 u_cpu.rf_ram.memory\[36\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08744_ u_cpu.rf_ram.memory\[136\]\[6\] _03782_ _03787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05956_ _01572_ _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06026__S1 _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08675_ _03680_ _03735_ _03742_ _00540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05887_ u_arbiter.i_wb_cpu_dbus_adr\[18\] _01512_ _01518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06726__I0 u_cpu.rf_ram.memory\[76\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08340__A2 _03526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07626_ _02751_ _03070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07557_ _02987_ _03022_ _03025_ _00139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_41_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06508_ _01638_ _02122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_10_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11526__CLK net432 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07488_ u_cpu.rf_ram.memory\[45\]\[5\] _02973_ _02977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06439_ u_cpu.rf_ram.memory\[136\]\[2\] u_cpu.rf_ram.memory\[137\]\[2\] u_cpu.rf_ram.memory\[138\]\[2\]
+ u_cpu.rf_ram.memory\[139\]\[2\] _01814_ _01942_ _02054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09227_ u_cpu.rf_ram.memory\[92\]\[4\] _04097_ _04100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07851__A1 _03193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09169__I _04057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09158_ _03980_ _04045_ _04051_ _00714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10738__A1 _05146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08109_ _03342_ _03382_ _03387_ _00329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06406__A2 _02020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11676__CLK net288 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09089_ u_cpu.rf_ram.memory\[37\]\[2\] _04007_ _04008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11120_ u_cpu.cpu.ctrl.i_iscomp _04467_ _05442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09356__A1 _04152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11051_ _05352_ _05392_ _05395_ _01264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11163__A1 _05454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10002_ _03115_ u_arbiter.i_wb_cpu_rdt\[29\] _04697_ _04698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_76_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07906__A2 _03255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05917__A1 _01537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10910__A1 _05278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09659__A2 _04384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11953_ _00649_ net440 u_cpu.rf_ram.memory\[126\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06717__I0 u_cpu.rf_ram.memory\[84\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12301__CLK net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08331__A2 _03529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10904_ u_cpu.rf_ram.memory\[84\]\[1\] _05303_ _05305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08248__I _03472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06342__A1 _01580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11884_ _00580_ net468 u_cpu.rf_ram.memory\[134\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10835_ u_cpu.rf_ram.memory\[83\]\[1\] _05258_ _05260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08095__A1 u_cpu.rf_ram.memory\[29\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10766_ _04832_ _05217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_40_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[60\] u_scanchain_local.module_data_in\[59\] net554 u_arbiter.o_wb_cpu_adr\[22\]
+ net22 u_scanchain_local.module_data_in\[60\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
X_12505_ _01184_ net168 u_cpu.rf_ram.memory\[83\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07842__A1 _03179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08890__I0 _03572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10697_ u_cpu.rf_ram.memory\[103\]\[6\] _05168_ _05173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12436_ _01115_ net160 u_cpu.rf_ram.memory\[101\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12367_ _01046_ net210 u_cpu.rf_ram.memory\[93\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11318_ _05562_ _01364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06799__I3 u_cpu.rf_ram.memory\[95\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12298_ _00980_ net94 u_cpu.rf_ram.memory\[30\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09347__A1 _04140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11249_ _05462_ _05512_ _05521_ _01336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09898__A2 _04453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout384_I net385 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06256__S1 _01676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05810_ _01455_ _01456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08570__A2 _03674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06790_ _02014_ _02400_ _02401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05741_ _01391_ _01368_ _01392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_fanout551_I net565 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10688__I _05163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08322__A2 _03514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08460_ u_cpu.rf_ram.memory\[141\]\[1\] _03610_ _03612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11549__CLK net339 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07411_ u_cpu.rf_ram.memory\[78\]\[1\] _02926_ _02928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08391_ _02857_ _03566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07997__I _03311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07342_ _02784_ _02875_ _02876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_50_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10968__A1 _05278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09822__A2 _04457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07833__A1 _03195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07273_ u_cpu.rf_ram.memory\[18\]\[5\] _02822_ _02826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09012_ _02981_ _03181_ _03957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06224_ _01570_ _01839_ _01840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06155_ _01702_ _01772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09717__I _04441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06086_ _01702_ _01703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09338__A1 _04154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09914_ _04607_ _04618_ _04619_ _04620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_63_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11145__A1 _05458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08010__A1 _02723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09845_ _04522_ _04561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09776_ _04498_ _04499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06988_ _01411_ _02593_ _02594_ _01374_ _02595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__05980__I _01596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08727_ _03763_ _03767_ _03776_ _00558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05939_ u_cpu.cpu.ctrl.o_ibus_adr\[30\] _01557_ _01558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07116__A3 _02701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09510__A1 u_cpu.rf_ram.memory\[33\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08313__A2 _03517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08658_ u_cpu.rf_ram.memory\[138\]\[7\] _03721_ _03732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10120__A2 _04619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12474__CLK net182 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07609_ u_cpu.rf_ram.memory\[48\]\[6\] _03052_ _03057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06875__A2 _02484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08589_ u_cpu.rf_ram.memory\[70\]\[2\] _03691_ _03692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10620_ u_arbiter.i_wb_cpu_rdt\[26\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[10\]
+ _05123_ _05124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08077__A1 _03353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10551_ _02890_ _04959_ _05083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07824__A1 _03186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06183__S0 _01798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10482_ _02787_ _05006_ _05037_ _05038_ _01052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06316__I _01627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12221_ _00904_ net350 u_cpu.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08624__I0 _03560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07348__S _02879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12152_ _00835_ net398 u_cpu.rf_ram.memory\[116\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06486__S1 _02099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11103_ _05428_ _05418_ _05429_ _02577_ _01282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09329__A1 _04145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12083_ _00766_ net448 u_cpu.rf_ram.memory\[120\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11136__A1 _05451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11034_ _05354_ _05380_ _05385_ _01257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06051__I _01667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08001__A1 _03262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09790__C _04511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08552__A2 _03656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11936_ _00632_ net462 u_cpu.rf_ram.memory\[128\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10111__A2 _04750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11867_ _00563_ net519 u_cpu.rf_ram.memory\[136\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08068__A1 u_cpu.rf_ram.memory\[64\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10818_ u_cpu.rf_ram.memory\[107\]\[2\] _05249_ _05250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09804__A2 _04457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11798_ _00494_ net368 u_cpu.rf_ram.memory\[73\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06618__A2 _02230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07815__A1 _03199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout132_I net157 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10749_ _05204_ _05201_ _05205_ _01152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11991__CLK net257 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07291__A2 _02833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12419_ _01098_ net357 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10178__A2 _04837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08240__A1 _03417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12347__CLK net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07960_ _03293_ _00274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06911_ u_cpu.rf_ram.memory\[128\]\[7\] u_cpu.rf_ram.memory\[129\]\[7\] u_cpu.rf_ram.memory\[130\]\[7\]
+ u_cpu.rf_ram.memory\[131\]\[7\] _01614_ _01616_ _02521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07891_ u_cpu.rf_ram.memory\[74\]\[4\] _03245_ _03248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09630_ u_arbiter.i_wb_cpu_dbus_dat\[26\] _04370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09740__A1 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08543__A2 _03659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06842_ _02081_ _02451_ _01603_ _02452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11371__CLK net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06554__A1 _01400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12497__CLK net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09561_ _04321_ _04322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06773_ u_cpu.rf_ram.memory\[36\]\[6\] u_cpu.rf_ram.memory\[37\]\[6\] u_cpu.rf_ram.memory\[38\]\[6\]
+ u_cpu.rf_ram.memory\[39\]\[6\] _01716_ _02109_ _02384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09205__C _02559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05724_ _01374_ _01375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08512_ _03641_ _00478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout45_I net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09492_ u_cpu.rf_ram.memory\[116\]\[6\] _04262_ _04267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07354__I0 _02864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08443_ _03500_ _03600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_24_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06401__S1 _01737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08374_ _03498_ _03549_ _03555_ _00426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07325_ u_cpu.rf_ram_if.wdata0_r\[4\] u_cpu.rf_ram_if.wdata1_r\[4\] _02844_ _02863_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_17_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06609__A2 _02221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07806__A1 _03193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06136__I _01706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07256_ _02773_ _02807_ _02815_ _00048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07282__A2 _02831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09559__A1 u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06207_ _01819_ _01822_ _01823_ _01824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07187_ _02733_ _02763_ _02764_ _00030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05975__I _01576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10169__A2 _04840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10413__I0 _04192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06138_ _01662_ _01755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07034__A2 _02586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08231__A1 _03405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06468__S1 _01968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08782__A2 _03806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06069_ _01685_ _01686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__11118__A1 u_cpu.cpu.genblk3.csr.mstatus_mie vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout410 net412 net410 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_120_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout421 net423 net421 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__11714__CLK net450 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout432 net433 net432 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_28_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout443 net444 net443 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout454 net455 net454 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_63_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout465 net467 net465 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_47_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09731__A1 _04450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout476 net538 net476 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_101_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09828_ _04470_ _04545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout487 net489 net487 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout498 net499 net498 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_115_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06739__C _01405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09759_ _02680_ _04482_ _04483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08298__A1 _03507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11721_ _00425_ net452 u_cpu.rf_ram.memory\[52\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11652_ _00356_ net220 u_cpu.rf_ram.memory\[60\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout50 net73 net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__07430__I _02939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout61 net62 net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_10603_ _05114_ _01097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout72 net73 net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_128_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout83 net84 net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_11583_ _00287_ net245 u_cpu.rf_ram.memory\[67\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout94 net95 net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_70_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08470__A1 _03602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10534_ u_cpu.rf_ram.memory\[95\]\[0\] _05073_ _05074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06046__I _01662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07273__A2 _02822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09785__C _04492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10791__I _05231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10465_ _04518_ _04434_ _05024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_6_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12204_ _00887_ net362 u_arbiter.i_wb_cpu_dbus_we vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_89_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10396_ _04977_ _01027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[23\] u_arbiter.i_wb_cpu_rdt\[20\] net541 u_arbiter.i_wb_cpu_dbus_dat\[17\]
+ net10 u_arbiter.i_wb_cpu_rdt\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
X_12135_ _00818_ net436 u_cpu.rf_ram.memory\[122\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08773__A2 _03803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06623__I2 u_cpu.rf_ram.memory\[94\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11394__CLK net297 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12066_ _00749_ net282 u_cpu.rf_ram.memory\[34\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08525__A2 _03647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11017_ u_cpu.rf_ram.memory\[86\]\[4\] _05372_ _05375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11127__I _05445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08289__A1 u_cpu.rf_ram.memory\[56\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11919_ _00615_ net144 u_cpu.rf_ram.memory\[12\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout347_I net349 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08436__I _03493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout514_I net515 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06147__S0 _01762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07110_ _02610_ _02611_ _02698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08090_ _03345_ _03369_ _03375_ _00322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08461__A1 _03593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07264__A2 _02819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06698__S1 _01693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07041_ u_cpu.rf_ram_if.rtrig1 _02646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10407__S _04983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05795__I _01441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07016__A2 _02616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11737__CLK net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10206__I _02690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09961__A1 _04528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08764__A2 _03794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08992_ _02966_ _03181_ _03945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10571__A2 _04467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07943_ _03266_ _03275_ _03282_ _00268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06870__S1 _01660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09713__A1 _04437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08516__A2 _03644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07874_ _03195_ _03230_ _03237_ _00244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06527__A1 _01423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07515__I _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09613_ _04294_ _04359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_95_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06825_ u_cpu.rf_ram.memory\[132\]\[6\] u_cpu.rf_ram.memory\[133\]\[6\] u_cpu.rf_ram.memory\[134\]\[6\]
+ u_cpu.rf_ram.memory\[135\]\[6\] _02061_ _02174_ _02436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_3_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09544_ u_arbiter.i_wb_cpu_dbus_dat\[2\] _04299_ _04307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06756_ _01590_ _02366_ _02367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07327__I0 _02864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09475_ _04255_ _04240_ _04256_ _00827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06687_ u_cpu.rf_ram.memory\[32\]\[5\] u_cpu.rf_ram.memory\[33\]\[5\] u_cpu.rf_ram.memory\[34\]\[5\]
+ u_cpu.rf_ram.memory\[35\]\[5\] _01767_ _01994_ _02299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08426_ _03587_ _00446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08357_ u_cpu.rf_ram.memory\[53\]\[5\] _03541_ _03545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12512__CLK net203 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09378__S _04186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07308_ _02849_ _02850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_71_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07255__A2 _02810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08288_ _03500_ _03501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07239_ _02731_ _02804_ _02805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09177__I _04057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10250_ _02689_ _03123_ _04885_ _04886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_106_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12662__CLK net159 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08204__A1 _03419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10181_ u_cpu.cpu.alu.cmp_r _02699_ _04847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xfanout240 net247 net240 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__06861__S1 _02109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout251 net254 net251 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__09704__A1 _04421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout262 net266 net262 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout273 net274 net273 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_115_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout284 net285 net284 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_134_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout295 net298 net295 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06613__S1 _01737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11704_ _00408_ net421 u_cpu.rf_ram.memory\[54\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12684_ u_cpu.rf_ram_if.wdata0_r\[1\] net232 u_cpu.rf_ram_if.wdata0_r\[0\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08691__A1 u_cpu.rf_ram.memory\[137\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[33\]_CLK net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12192__CLK net498 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11635_ _00339_ net175 u_cpu.rf_ram.memory\[62\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09640__B1 _04295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11566_ _00270_ net341 u_cpu.rf_ram.memory\[75\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10517_ _05044_ _05060_ _05063_ _01062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11497_ _00201_ net178 u_cpu.rf_ram.memory\[17\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_u_scanchain_local.scan_flop\[48\]_CLK net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10448_ _04566_ _04503_ _04602_ _05008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10002__A1 _03115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09943__A1 _04601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08746__A2 _03777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10379_ u_cpu.rf_ram.memory\[109\]\[4\] _04965_ _04968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12118_ _00801_ net127 u_cpu.rf_ram.memory\[11\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10470__B _05025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06852__S1 _01633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout297_I net298 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12049_ _00732_ net271 u_cpu.rf_ram.memory\[92\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09171__A2 _04059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06604__S1 _01717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07182__A1 _02748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06610_ u_cpu.rf_ram.memory\[96\]\[4\] u_cpu.rf_ram.memory\[97\]\[4\] u_cpu.rf_ram.memory\[98\]\[4\]
+ u_cpu.rf_ram.memory\[99\]\[4\] _02125_ _01693_ _02223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_111_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07590_ _02998_ _03037_ _03045_ _00152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09550__I _04311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10069__A1 _04490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06541_ _02144_ _02146_ _02149_ _02154_ _01925_ _02155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_46_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06368__S0 _01871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09260_ u_cpu.rf_ram.memory\[34\]\[1\] _04118_ _04120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06472_ _01630_ _02085_ _02086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07485__A2 _02969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08211_ _02846_ u_cpu.rf_ram.memory\[5\]\[0\] _03451_ _03452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09191_ _04072_ _04059_ _04073_ _00725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08142_ _03406_ _03407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12685__CLK net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08073_ _03349_ _03357_ _03364_ _00316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08985__A2 _03934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07024_ u_cpu.cpu.mem_bytecnt\[1\] _02628_ _02629_ _02630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10792__A2 _05233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06414__I _01704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08737__A2 _03778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10544__A2 _05072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06599__I1 u_cpu.rf_ram.memory\[33\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06843__S1 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08975_ u_cpu.rf_ram.memory\[126\]\[0\] _03935_ _03936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07926_ _03270_ _03255_ _03271_ _00262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12065__CLK net284 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07012__I2 u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07857_ _03199_ _03217_ _03226_ _00238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10600__S _05111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06808_ u_cpu.rf_ram.memory\[64\]\[6\] u_cpu.rf_ram.memory\[65\]\[6\] u_cpu.rf_ram.memory\[66\]\[6\]
+ u_cpu.rf_ram.memory\[67\]\[6\] _01798_ _02040_ _02419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_28_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07788_ _03180_ _03181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_45_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09527_ net8 _01450_ _04292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_77_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06739_ _02344_ _02346_ _02348_ _02350_ _01405_ _02351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_24_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06359__S0 _01640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09458_ _04238_ _04245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08673__A1 _03678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11902__CLK net459 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10480__A1 _04516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08409_ _03285_ _03062_ _03578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_71_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09389_ _03870_ _03034_ _04202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_40_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11420_ _00124_ net297 u_cpu.rf_ram.memory\[44\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07228__A2 _02792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09622__B1 _04359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08976__A2 _03934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11351_ _00055_ net69 u_cpu.rf_ram.memory\[18\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06987__A1 _01408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06531__S0 _02029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10783__A2 _05224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10302_ u_cpu.cpu.ctrl.o_ibus_adr\[7\] _04915_ _04917_ u_cpu.cpu.ctrl.o_ibus_adr\[8\]
+ _04920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11282_ u_cpu.rf_ram.memory\[89\]\[4\] _05539_ _05542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08728__A2 _03698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10233_ u_arbiter.i_wb_cpu_dbus_adr\[25\] u_arbiter.i_wb_cpu_dbus_adr\[24\] _04873_
+ _04876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10535__A2 _05072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07356__S _02878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12408__CLK net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10164_ u_cpu.rf_ram.memory\[31\]\[0\] _04837_ _04838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07400__A2 _02714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06834__S1 _02071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10095_ u_cpu.cpu.immdec.imm19_12_20\[6\] _04772_ _04782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05962__A2 _01578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11432__CLK net368 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12558__CLK net212 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06211__I0 u_cpu.rf_ram.memory\[128\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08900__A2 _03882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06762__I1 u_cpu.rf_ram.memory\[49\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10997_ u_cpu.rf_ram.memory\[110\]\[5\] _05355_ _05362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11582__CLK net340 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08664__A1 _03666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10471__A1 _04510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10471__B2 _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12667_ _01346_ net287 u_cpu.rf_ram.memory\[89\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11618_ _00322_ net103 u_cpu.rf_ram.memory\[29\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12598_ _01277_ net279 u_cpu.rf_ram.memory\[88\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06662__C _01807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08967__A2 _03923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout212_I net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11549_ _00253_ net339 u_cpu.rf_ram.memory\[74\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11140__I _02762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10774__A2 _05221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09916__A1 _04484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12088__CLK net438 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06825__S1 _02174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08760_ u_cpu.rf_ram.memory\[135\]\[4\] _03794_ _03797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05972_ _01580_ _01586_ _01588_ _01589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07711_ net8 _01450_ _03132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08691_ u_cpu.rf_ram.memory\[137\]\[2\] _03753_ _03754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07642_ _03081_ _03065_ _03082_ _00167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11925__CLK net236 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07573_ _03018_ _03034_ _03035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09312_ u_cpu.rf_ram.memory\[120\]\[4\] _04148_ _04153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07014__B _02620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06524_ _01751_ _02137_ _01755_ _02138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08655__A1 _03680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09243_ u_cpu.rf_ram.memory\[35\]\[2\] _04109_ _04110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06455_ _01418_ _02069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06386_ _01638_ _02001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09174_ u_cpu.rf_ram.memory\[90\]\[1\] _04059_ _04062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06269__I0 u_cpu.rf_ram.memory\[32\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08958__A2 _03922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08125_ u_cpu.rf_ram.memory\[62\]\[1\] _03395_ _03397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09080__A1 _03988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06969__A1 _01394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06144__I _01648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08056_ u_cpu.rf_ram.memory\[65\]\[7\] _03336_ _03354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07630__A2 _03064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09907__A1 _04443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07007_ u_cpu.cpu.decode.opcode\[0\] _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_1_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10517__A2 _05060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11455__CLK net370 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11190__A2 _05476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08958_ _03900_ _03922_ _03925_ _00640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09391__S _04203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07909_ _03253_ _03260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08889_ _03877_ _00619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10920_ _05313_ _05314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_79_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10851_ _02981_ _05243_ _05269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08646__A1 _03671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10782_ _05211_ _05220_ _05227_ _01163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10453__A1 _04560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12521_ _01200_ net296 u_cpu.rf_ram.memory\[69\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06763__B _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12452_ _01131_ net87 u_cpu.rf_ram.memory\[103\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11403_ _00107_ net218 u_cpu.rf_ram.memory\[46\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12383_ _01062_ net195 u_cpu.rf_ram.memory\[94\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06504__S0 _02001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10756__A2 _05201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06054__I _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11334_ _00038_ net60 u_cpu.rf_ram.memory\[21\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07621__A2 _03064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11265_ _02909_ _05524_ _05531_ _01342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09365__I _04185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10216_ _04866_ _00958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11196_ _05444_ _05489_ _05491_ _01313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11181__A2 _05477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10147_ u_cpu.rf_ram.memory\[32\]\[4\] _04818_ _04825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11948__CLK net461 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09126__A2 _02563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10078_ _04753_ _04764_ _04765_ _04766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_47_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07613__I _02739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06735__I1 u_cpu.rf_ram.memory\[129\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10692__A1 _05140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout162_I net163 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06360__A2 _01974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10444__A1 _03118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10995__A2 _05349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06240_ _01630_ _01855_ _01856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09598__C1 _04327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06171_ _01575_ _01788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07612__A2 _03049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11478__CLK net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09930_ u_cpu.cpu.immdec.imm24_20\[1\] _04629_ _04633_ u_cpu.cpu.immdec.imm24_20\[2\]
+ _04634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_89_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10415__S _04983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09861_ _04525_ _04563_ _04576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05736__C _01386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09208__C _02676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06179__A2 _01794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11172__A2 _03020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08812_ u_cpu.rf_ram.memory\[133\]\[6\] _03822_ _03831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09792_ _04513_ _00887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_86_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05926__A2 u_cpu.cpu.ctrl.o_ibus_adr\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09117__A2 _04019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08743_ _03759_ _03779_ _03786_ _00564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05955_ _01571_ _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07128__A1 _02535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08876__A1 _03832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08674_ u_cpu.rf_ram.memory\[39\]\[5\] _03738_ _03742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05886_ u_cpu.cpu.ctrl.o_ibus_adr\[17\] _01511_ u_cpu.cpu.ctrl.o_ibus_adr\[18\] _01517_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_81_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07625_ _03068_ _03064_ _03069_ _00163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07556_ u_cpu.rf_ram.memory\[41\]\[1\] _03023_ _03025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09676__I0 u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06507_ _02004_ _02120_ _01723_ _02121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_42_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07300__A1 u_cpu.rf_ram.memory\[20\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07487_ _02907_ _02969_ _02976_ _00118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05978__I _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09226_ _04066_ _04093_ _04099_ _00735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12253__CLK net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06438_ _02025_ _02052_ _01810_ _02053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09157_ u_cpu.rf_ram.memory\[91\]\[3\] _04049_ _04051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06369_ _01672_ _01983_ _01873_ _01984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_33_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08108_ u_cpu.rf_ram.memory\[63\]\[2\] _03386_ _03387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09088_ _04002_ _04007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07603__A2 _03052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08039_ _03070_ _03342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_104_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09356__A2 _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11050_ u_cpu.rf_ram.memory\[87\]\[1\] _05393_ _05395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06009__I3 u_cpu.rf_ram.memory\[19\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10001_ _01443_ u_arbiter.i_wb_cpu_rdt\[13\] _04697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_77_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05917__A2 _01535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10910__A2 _05302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06758__B _01588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11952_ _00648_ net453 u_cpu.rf_ram.memory\[126\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10903_ _05268_ _05302_ _05304_ _01207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11883_ _00579_ net518 u_cpu.rf_ram.memory\[134\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06342__A2 _01956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08619__A1 _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10834_ _05199_ _05257_ _05259_ _01183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06049__I _01665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09292__A1 _04072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10765_ _05215_ _05202_ _05216_ _01157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12504_ _01183_ net185 u_cpu.rf_ram.memory\[83\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10696_ _05144_ _05165_ _05172_ _01132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06496__I3 u_cpu.rf_ram.memory\[39\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11226__I0 _02869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[53\] u_scanchain_local.module_data_in\[52\] net561 u_arbiter.o_wb_cpu_adr\[15\]
+ net29 u_scanchain_local.module_data_in\[53\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_12_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12435_ _01114_ net160 u_cpu.rf_ram.memory\[101\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09044__A1 u_cpu.rf_ram.memory\[123\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11620__CLK net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12366_ _01045_ net210 u_cpu.rf_ram.memory\[93\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11317_ _04032_ u_cpu.rf_ram_if.rreq_r _05562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_99_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12297_ _00979_ net103 u_cpu.rf_ram.memory\[30\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11770__CLK net490 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09347__A2 _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11248_ u_cpu.rf_ram.memory\[98\]\[7\] _05510_ _05521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06405__I0 u_cpu.rf_ram.memory\[112\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11179_ _05476_ _05481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout377_I net381 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12126__CLK net405 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05740_ u_cpu.cpu.csr_imm _01391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_23_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07343__I _02876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10665__A1 u_cpu.rf_ram.memory\[102\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout544_I net546 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06333__A2 _01948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07410_ _02889_ _02925_ _02927_ _00090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12276__CLK net533 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08390_ _03565_ _00432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07341_ _02719_ _02781_ _02875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__10968__A2 _05336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11090__A1 _01386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07272_ _02763_ _02818_ _02825_ _00054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07833__A2 _03205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05844__A1 u_arbiter.i_wb_cpu_dbus_adr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09011_ _03919_ _03947_ _03956_ _00662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06223_ u_cpu.rf_ram.memory\[8\]\[1\] u_cpu.rf_ram.memory\[9\]\[1\] u_cpu.rf_ram.memory\[10\]\[1\]
+ u_cpu.rf_ram.memory\[11\]\[1\] _01574_ _01838_ _01839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_121_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06154_ _01766_ _01769_ _01770_ _01771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_144_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07597__A1 _02980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06085_ _01567_ _01702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07518__I _02912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09913_ _04528_ _04610_ _04459_ _04619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_99_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09844_ _04444_ _04560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08010__A2 _02923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09775_ _04464_ _04493_ _04498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06987_ _01408_ _01371_ _02594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_101_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08726_ u_cpu.rf_ram.memory\[49\]\[7\] _03765_ _03776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05938_ u_cpu.cpu.ctrl.o_ibus_adr\[29\] u_cpu.cpu.ctrl.o_ibus_adr\[28\] u_cpu.cpu.ctrl.o_ibus_adr\[27\]
+ _01548_ _01557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_27_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06297__C _01757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10656__A1 _05146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08657_ _03682_ _03723_ _03731_ _00533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05869_ _01502_ _01499_ _01503_ _01504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06324__A2 _01926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10120__A3 _04801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07608_ _02996_ _03049_ _03056_ _00159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08588_ _03686_ _03691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_74_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07539_ _02992_ _03007_ _03013_ _00133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09274__A1 _04074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11643__CLK net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06707__S0 _02136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11081__A1 u_cpu.rf_ram.memory\[88\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10550_ _05057_ _05073_ _05082_ _01076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06183__S1 _01799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09209_ _04078_ _04088_ _00729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10481_ u_cpu.cpu.immdec.imm30_25\[0\] _04630_ _05006_ _05038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_87_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12220_ _00903_ net353 u_cpu.cpu.decode.op26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11793__CLK net352 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07588__A1 _02996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12151_ _00834_ net401 u_cpu.rf_ram.memory\[116\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07428__I _02937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11102_ _01382_ _01393_ _05417_ _05429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_81_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09329__A2 _04161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12082_ _00765_ net436 u_cpu.rf_ram.memory\[120\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11033_ u_cpu.rf_ram.memory\[111\]\[2\] _05384_ _05385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08001__A2 _03312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06012__A1 _01619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10895__A1 _05284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12299__CLK net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09501__A2 _04271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10647__A1 _05140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11935_ _00631_ net454 u_cpu.rf_ram.memory\[128\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11866_ _00562_ net518 u_cpu.rf_ram.memory\[136\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10817_ _05244_ _05249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_18_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11797_ _00493_ net371 u_cpu.rf_ram.memory\[73\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06079__A1 _01691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10748_ u_cpu.rf_ram.memory\[79\]\[1\] _05202_ _05205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05826__A1 _01434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout125_I net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10679_ _05148_ _05152_ _05161_ _01126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_12418_ _01097_ net264 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07579__A1 _02987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12349_ _01028_ net125 u_cpu.rf_ram.memory\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08240__A2 _03461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07338__I _02872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout494_I net507 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06910_ _01830_ _02519_ _01628_ _02520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07890_ _03191_ _03241_ _03247_ _00250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11516__CLK net400 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09740__A2 _01433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06841_ u_cpu.rf_ram.memory\[16\]\[7\] u_cpu.rf_ram.memory\[17\]\[7\] u_cpu.rf_ram.memory\[18\]\[7\]
+ u_cpu.rf_ram.memory\[19\]\[7\] _01598_ _01599_ _02451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_116_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06554__A2 _02167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09560_ _04294_ _04321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_7_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06772_ _01988_ _02382_ _02107_ _02383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_36_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08511_ _03576_ u_cpu.rf_ram.memory\[13\]\[7\] _03632_ _03641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05723_ u_cpu.cpu.decode.opcode\[2\] _01374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09491_ _04251_ _04259_ _04266_ _00833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07503__A1 u_cpu.rf_ram.memory\[44\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11666__CLK net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08442_ _03598_ _03590_ _03599_ _00450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout38_I net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07801__I _03074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08373_ u_cpu.rf_ram.memory\[52\]\[3\] _03553_ _03555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07324_ _02862_ _00069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11063__A1 u_cpu.rf_ram.memory\[87\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10810__A1 _03033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09008__A1 u_cpu.rf_ram.memory\[125\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07255_ u_cpu.rf_ram.memory\[81\]\[6\] _02810_ _02815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06206_ _01602_ _01823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07186_ u_cpu.rf_ram.memory\[82\]\[4\] _02753_ _02764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06617__I0 u_cpu.rf_ram.memory\[112\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06137_ u_cpu.rf_ram.memory\[116\]\[0\] u_cpu.rf_ram.memory\[117\]\[0\] u_cpu.rf_ram.memory\[118\]\[0\]
+ u_cpu.rf_ram.memory\[119\]\[0\] _01752_ _01753_ _01754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08231__A2 _03461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06068_ _01581_ _01685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout400 net402 net400 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout411 net412 net411 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_87_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07990__A1 _03272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout422 net423 net422 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_134_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout433 net434 net433 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_58_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10326__B1 _04931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout444 net447 net444 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_63_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout455 net460 net455 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout466 net467 net466 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_63_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09827_ _04412_ _04434_ _04453_ _04427_ _04486_ _04544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
Xfanout477 net484 net477 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_24_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10877__A1 _05286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09731__A2 _04453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout488 net489 net488 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XTAP_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout499 net506 net499 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_86_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06545__A2 _02158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06396__I2 u_cpu.rf_ram.memory\[98\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09758_ _04481_ _04482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08709_ _03765_ _03766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09689_ _04413_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[0\] _04414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09495__A1 _04255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08298__A2 _03488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11720_ _00424_ net418 u_cpu.rf_ram.memory\[52\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11651_ _00355_ net216 u_cpu.rf_ram.memory\[60\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout40 net42 net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_80_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout51 net55 net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_126_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10602_ u_arbiter.i_wb_cpu_rdt\[18\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[2\]
+ _05111_ _05114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11054__A1 _05354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout62 net72 net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_11582_ _00286_ net340 u_cpu.rf_ram.memory\[68\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout73 net109 net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_141_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout84 net92 net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout95 net97 net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_80_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10801__A1 u_cpu.rf_ram.memory\[106\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10533_ _05071_ _05073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_7_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08470__A2 _03610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10464_ _02701_ _04630_ _05022_ _05023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12203_ _00886_ net384 u_cpu.cpu.decode.opcode\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10395_ _04192_ u_cpu.rf_ram.memory\[3\]\[3\] _04973_ _04977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_48_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07158__I _02739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11539__CLK net242 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12134_ _00817_ net438 u_cpu.rf_ram.memory\[122\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06062__I _01678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06623__I3 u_cpu.rf_ram.memory\[95\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[16\] u_arbiter.i_wb_cpu_rdt\[13\] net542 u_arbiter.i_wb_cpu_dbus_dat\[10\]
+ net11 u_arbiter.i_wb_cpu_rdt\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
X_12065_ _00748_ net284 u_cpu.rf_ram.memory\[34\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10868__A1 _05280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11016_ _05357_ _05368_ _05374_ _01250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07733__A1 _03071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06387__I2 u_cpu.rf_ram.memory\[110\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08289__A2 _03495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10096__A2 _04780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11918_ _00614_ net457 u_cpu.rf_ram.memory\[130\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11849_ _00545_ net508 u_cpu.rf_ram.memory\[137\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout242_I net246 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11143__I _02767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11045__A1 _05300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06147__S1 _01763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08461__A2 _03609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout507_I net537 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07040_ _02645_ u_cpu.cpu.o_wdata0 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06472__A1 _01630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08452__I _03509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07016__A3 _00728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07068__I _01401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06224__A1 _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09961__A2 _04567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08991_ _03919_ _03935_ _03944_ _00654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07972__A1 u_cpu.rf_ram.memory\[68\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07942_ u_cpu.rf_ram.memory\[75\]\[5\] _03278_ _03282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09713__A2 _04418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07873_ u_cpu.rf_ram.memory\[77\]\[5\] _03233_ _03237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06527__A2 _02128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09612_ u_arbiter.i_wb_cpu_dbus_dat\[20\] _04352_ _04358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06824_ _01611_ _02434_ _02435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07017__B _02575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09543_ _04285_ _04305_ _04306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06755_ u_cpu.rf_ram.memory\[28\]\[6\] u_cpu.rf_ram.memory\[29\]\[6\] u_cpu.rf_ram.memory\[30\]\[6\]
+ u_cpu.rf_ram.memory\[31\]\[6\] _02084_ _01577_ _02366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_77_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11284__A1 u_cpu.rf_ram.memory\[89\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09474_ u_cpu.rf_ram.memory\[115\]\[7\] _04238_ _04256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_u_scanchain_local.scan_flop\[64\]_SE net554 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06686_ _01882_ _02297_ _02298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08425_ _03576_ u_cpu.rf_ram.memory\[15\]\[7\] _03578_ _03587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_52_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09229__A1 u_cpu.rf_ram.memory\[92\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11036__A1 _05357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08356_ _03501_ _03537_ _03544_ _00419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07307_ _02726_ _02578_ _02788_ _02848_ _02849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_50_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08287_ _02761_ _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06302__I2 u_cpu.rf_ram.memory\[90\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05986__I _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07238_ _02803_ _02804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_30_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07169_ _02748_ u_cpu.rf_ram_if.wdata1_r\[2\] _02749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08204__A2 _03440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10180_ _04833_ _04837_ _04846_ _00942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11831__CLK net478 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout230 net231 net230 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout241 net246 net241 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_43_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09704__A2 _04423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout252 net253 net252 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_75_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout263 net264 net263 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_86_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout274 net275 net274 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_74_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout285 net289 net285 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__06518__A2 _02131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout296 net297 net296 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_21_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10132__I _02744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11981__CLK net410 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11703_ _00407_ net330 u_cpu.rf_ram.memory\[54\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12683_ _01361_ net496 u_cpu.cpu.state.ibus_cyc vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12337__CLK net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08691__A2 _03753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06057__I _01673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11634_ _00338_ net175 u_cpu.rf_ram.memory\[62\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11565_ _00269_ net341 u_cpu.rf_ram.memory\[75\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09640__A1 u_arbiter.i_wb_cpu_rdt\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09640__B2 u_arbiter.i_wb_cpu_dbus_dat\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05896__I _01455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09368__I _02854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10516_ u_cpu.rf_ram.memory\[94\]\[1\] _05061_ _05063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12487__CLK net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11361__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10250__A2 _03123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11496_ _00200_ net140 u_cpu.rf_ram.memory\[17\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10447_ _02535_ _05006_ _05007_ _04732_ _01048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10389__I0 _04184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10002__A2 u_arbiter.i_wb_cpu_rdt\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09943__A2 _04609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10378_ _04821_ _04961_ _04967_ _01019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12117_ _00800_ net128 u_cpu.rf_ram.memory\[11\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10243__S _04848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10470__C _04582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07616__I _03061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12048_ _00731_ net379 u_cpu.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout192_I net193 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07182__A2 u_cpu.rf_ram_if.wdata1_r\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10977__I _02739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout457_I net459 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06540_ _02150_ _02152_ _02153_ _02154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_34_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08131__A1 _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06368__S1 _01676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06471_ u_cpu.rf_ram.memory\[28\]\[3\] u_cpu.rf_ram.memory\[29\]\[3\] u_cpu.rf_ram.memory\[30\]\[3\]
+ u_cpu.rf_ram.memory\[31\]\[3\] _02084_ _01634_ _02085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_34_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08210_ _03450_ _03451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__11018__A1 _05359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06693__A1 _02117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09190_ u_cpu.rf_ram.memory\[90\]\[6\] _04064_ _04073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11704__CLK net421 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08141_ _02966_ _03005_ _03406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08434__A2 _03591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08072_ u_cpu.rf_ram.memory\[64\]\[5\] _03360_ _03364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06996__A2 _02602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07023_ _02532_ _02624_ _02629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10217__I _02690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11854__CLK net510 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08198__A1 _03412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09934__A2 _04627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07945__A1 _03268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08974_ _03933_ _03935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07925_ u_cpu.rf_ram.memory\[76\]\[7\] _03253_ _03271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09698__A1 _03114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07856_ u_cpu.rf_ram.memory\[139\]\[7\] _03215_ _03226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07012__I3 u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06807_ _02411_ _02413_ _02415_ _02417_ _01757_ _02418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_42_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07787_ _02729_ _03003_ _03180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09526_ net36 _04289_ _04290_ _04291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06738_ _02060_ _02349_ _01644_ _02350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07261__I _02817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06359__S1 _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09457_ _03902_ _04244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06669_ u_cpu.rf_ram.memory\[24\]\[5\] u_cpu.rf_ram.memory\[25\]\[5\] u_cpu.rf_ram.memory\[26\]\[5\]
+ u_cpu.rf_ram.memory\[27\]\[5\] _01622_ _01625_ _02281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_52_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08673__A2 _03734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06523__I2 u_cpu.rf_ram.memory\[118\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08408_ _03577_ _00438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11009__A1 _05347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11384__CLK net217 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10480__A2 _04650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09388_ _04201_ _00795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08339_ u_cpu.rf_ram.memory\[54\]\[6\] _03529_ _03534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09622__A1 u_arbiter.i_wb_cpu_rdt\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11350_ _00054_ net67 u_cpu.rf_ram.memory\[18\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06987__A2 _01371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10301_ _04919_ _00990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06531__S1 _01768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11281_ _02903_ _05535_ _05541_ _01348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_4_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08189__A1 _03367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10232_ _04875_ _00965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06295__S0 _01752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10163_ _04835_ _04837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_48_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10094_ u_cpu.cpu.immdec.imm19_12_20\[7\] _04572_ _04781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[9\] u_arbiter.i_wb_cpu_rdt\[6\] net544 u_arbiter.i_wb_cpu_dbus_dat\[3\]
+ net12 u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_43_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06211__I1 u_cpu.rf_ram.memory\[129\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06762__I2 u_cpu.rf_ram.memory\[50\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08267__I _02738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11727__CLK net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10996_ _02767_ _05361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07171__I _02750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08113__A1 _03347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09861__A1 _04525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08664__A2 _03734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10471__A2 _04560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12666_ _01345_ net286 u_cpu.rf_ram.memory\[89\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11617_ _00321_ net103 u_cpu.rf_ram.memory\[29\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11877__CLK net516 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12597_ _01276_ net279 u_cpu.rf_ram.memory\[88\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07120__B _02704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11548_ _00252_ net339 u_cpu.rf_ram.memory\[74\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout205_I net207 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11479_ _00183_ net122 u_cpu.rf_ram.memory\[4\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08730__I _03777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06286__S0 _01736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05971_ _01587_ _01588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07710_ _01409_ _02559_ _03130_ _03131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__12502__CLK net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08690_ _03746_ _03753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09561__I _04321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07155__A2 _02736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08352__A1 _03494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07641_ u_cpu.rf_ram.memory\[47\]\[5\] _03072_ _03082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11743__D _00000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06753__I2 u_cpu.rf_ram.memory\[18\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11239__A1 _05451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07572_ _03033_ _03034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05961__I0 u_cpu.rf_ram.memory\[8\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08104__A1 _03335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09311_ _03909_ _04152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_62_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06523_ u_cpu.rf_ram.memory\[116\]\[3\] u_cpu.rf_ram.memory\[117\]\[3\] u_cpu.rf_ram.memory\[118\]\[3\]
+ u_cpu.rf_ram.memory\[119\]\[3\] _02136_ _01753_ _02137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_34_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09852__A1 _04475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09242_ _04104_ _04109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_61_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06454_ u_cpu.rf_ram.memory\[12\]\[3\] u_cpu.rf_ram.memory\[13\]\[3\] u_cpu.rf_ram.memory\[14\]\[3\]
+ u_cpu.rf_ram.memory\[15\]\[3\] _01583_ _01841_ _02068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA_fanout20_I net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09173_ _03899_ _04061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06385_ _01566_ _01964_ _01976_ _01999_ _02000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_120_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08124_ _03335_ _03394_ _03396_ _00335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06425__I _01584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06969__A2 _02576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07091__A1 _02676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08055_ _03086_ _03353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07006_ _02532_ _02613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09907__A2 _04546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06277__S0 _01721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08591__A1 u_cpu.rf_ram.memory\[70\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07394__A2 _02901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06160__I _01397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08957_ u_cpu.rf_ram.memory\[127\]\[1\] _03923_ _03925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12182__CLK net389 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[32\]_CLK net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10611__S _05117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07908_ _03070_ _03259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08888_ _03570_ u_cpu.rf_ram.memory\[12\]\[4\] _03872_ _03877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09391__I0 _04184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08343__A1 _02786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07839_ _03215_ _03216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_17_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10850_ _04807_ _05268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_u_scanchain_local.scan_flop\[47\]_CLK net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09509_ _04249_ _04270_ _04277_ _00840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10781_ u_cpu.rf_ram.memory\[105\]\[4\] _05224_ _05227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12520_ _01199_ net296 u_cpu.rf_ram.memory\[69\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12451_ _01130_ net87 u_cpu.rf_ram.memory\[103\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11402_ _00106_ net217 u_cpu.rf_ram.memory\[46\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06409__B2 _02023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05880__A2 _01512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12382_ _01061_ net196 u_cpu.rf_ram.memory\[94\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09071__A2 _03995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06504__S1 _01717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11333_ _00037_ net59 u_cpu.rf_ram.memory\[21\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11264_ u_cpu.rf_ram.memory\[100\]\[5\] _05527_ _05531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10215_ u_arbiter.i_wb_cpu_dbus_adr\[17\] u_arbiter.i_wb_cpu_dbus_adr\[16\] _04861_
+ _04866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12525__CLK net345 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11195_ u_cpu.rf_ram.memory\[24\]\[0\] _05490_ _05491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10146_ _04823_ _04824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10077_ _04561_ _04502_ _04602_ _04765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08334__A1 _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09531__B1 _04295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09834__A1 _04545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout155_I net156 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10979_ _05348_ _05349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_44_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10444__A2 _05004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout322_I net323 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12649_ _01328_ net134 u_cpu.rf_ram.memory\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09598__B1 _04321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12055__CLK net271 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06170_ _01612_ _01787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_11_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10990__I _02757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09860_ _04552_ _04575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08573__A1 u_cpu.rf_ram.memory\[71\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08811_ _03506_ _03830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09791_ _02633_ _04482_ _04508_ _04512_ _04513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10380__A1 _04824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08742_ u_cpu.rf_ram.memory\[136\]\[5\] _03782_ _03786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05954_ u_cpu.raddr\[0\] _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout68_I net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07804__I _03077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08673_ _03678_ _03734_ _03741_ _00539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05885_ u_cpu.cpu.ctrl.o_ibus_adr\[18\] u_cpu.cpu.ctrl.o_ibus_adr\[17\] u_cpu.cpu.ctrl.o_ibus_adr\[16\]
+ _01508_ _01516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__06336__B1 _01949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08876__A2 _03860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07624_ u_cpu.rf_ram.memory\[47\]\[1\] _03065_ _03069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07555_ _02980_ _03022_ _03024_ _00138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_59_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09825__A1 _01409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09676__I1 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06864__B _01731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06506_ u_cpu.rf_ram.memory\[104\]\[3\] u_cpu.rf_ram.memory\[105\]\[3\] u_cpu.rf_ram.memory\[106\]\[3\]
+ u_cpu.rf_ram.memory\[107\]\[3\] _02005_ _01892_ _02120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_50_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07687__I0 _02873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07486_ u_cpu.rf_ram.memory\[45\]\[4\] _02973_ _02976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07300__A2 _02832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09225_ u_cpu.rf_ram.memory\[92\]\[3\] _04097_ _04099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06583__C _01784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06437_ _02026_ _02038_ _02051_ _02052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_33_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09156_ _03977_ _04045_ _04050_ _00713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06155__I _01702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06368_ u_cpu.rf_ram.memory\[56\]\[2\] u_cpu.rf_ram.memory\[57\]\[2\] u_cpu.rf_ram.memory\[58\]\[2\]
+ u_cpu.rf_ram.memory\[59\]\[2\] _01871_ _01676_ _01983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09053__A2 _03978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08107_ _03381_ _03386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11422__CLK net291 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10606__S _05111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07695__B _03116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06498__S0 _01705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09087_ _03975_ _04003_ _04006_ _00688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08800__A2 _03822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06299_ _01687_ _01915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05994__I _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08038_ _03340_ _03337_ _03341_ _00304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06811__A1 _01778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08370__I _03548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10000_ _04500_ _04687_ _04694_ _04696_ _00912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__08564__A1 u_cpu.rf_ram.memory\[71\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11572__CLK net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12698__CLK net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09989_ _01443_ u_arbiter.i_wb_cpu_rdt\[12\] _04686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__10371__A1 _04808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08316__A1 _03501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11951_ _00647_ net453 u_cpu.rf_ram.memory\[126\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08867__A2 _03863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10902_ u_cpu.rf_ram.memory\[84\]\[0\] _05303_ _05304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06878__A1 _01649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11882_ _00578_ net470 u_cpu.rf_ram.memory\[134\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10833_ u_cpu.rf_ram.memory\[83\]\[0\] _05258_ _05259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09816__A1 _04468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08619__A2 _03701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12078__CLK net319 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10764_ u_cpu.rf_ram.memory\[79\]\[6\] _05207_ _05216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12503_ _01182_ net41 u_cpu.rf_ram.memory\[107\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10695_ u_cpu.rf_ram.memory\[103\]\[5\] _05168_ _05172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12434_ _01113_ net87 u_cpu.rf_ram.memory\[101\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09044__A2 _03978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_scanchain_local.scan_flop\[46\] u_scanchain_local.module_data_in\[45\] net558 u_arbiter.o_wb_cpu_adr\[8\]
+ net26 u_scanchain_local.module_data_in\[46\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_86_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12365_ _01044_ net210 u_cpu.rf_ram.memory\[93\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11316_ _05561_ _01363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06802__A1 _01740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12296_ _00978_ net97 u_cpu.rf_ram.memory\[30\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11247_ _05460_ _05512_ _05520_ _01335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11178_ _05449_ _05477_ _05480_ _01306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10362__A1 _04953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10129_ _04809_ _04811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08307__A1 _03485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10114__A1 _02676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11146__I _02772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06869__A1 _02117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10665__A2 _05152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout537_I net538 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07340_ _02874_ _00073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11445__CLK net325 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07294__A1 u_cpu.rf_ram.memory\[20\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07271_ u_cpu.rf_ram.memory\[18\]\[4\] _02822_ _02825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06097__A2 _01608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09010_ u_cpu.rf_ram.memory\[125\]\[7\] _03945_ _03956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06222_ _01576_ _01838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_129_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05844__A2 _01453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06153_ _01418_ _01770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11595__CLK net251 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08794__A1 _03813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07597__A2 _03048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08190__I _03438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06084_ _01697_ _01700_ _01701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09912_ _04608_ _04548_ _04561_ _04601_ _04617_ _04618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_28_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08546__A1 _03600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09843_ u_arbiter.i_wb_cpu_rdt\[21\] u_arbiter.i_wb_cpu_rdt\[5\] _01447_ _04559_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09774_ _04426_ _04497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06986_ u_cpu.cpu.branch_op u_cpu.cpu.decode.opcode\[0\] _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05937_ _01489_ _01555_ _01556_ u_arbiter.o_wb_cpu_adr\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08725_ _03761_ _03767_ _03775_ _00557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_73_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08849__A2 _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08656_ u_cpu.rf_ram.memory\[138\]\[6\] _03726_ _03731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10656__A2 _05133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05868_ _01502_ _01499_ _01455_ _01503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__12220__CLK net353 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07607_ u_cpu.rf_ram.memory\[48\]\[5\] _03052_ _03056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08587_ _03671_ _03687_ _03690_ _00504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05799_ _01441_ _01446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_109_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05989__I _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08365__I _03548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07538_ u_cpu.rf_ram.memory\[51\]\[3\] _03011_ _03013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06707__S1 _01707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07285__A1 u_cpu.rf_ram.memory\[20\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07469_ u_cpu.rf_ram.memory\[46\]\[7\] _02953_ _02964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12370__CLK net359 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09397__S _04203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09208_ _02703_ _04087_ _00703_ _02676_ _04088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_10480_ _04516_ _04650_ _05036_ _05037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06883__I1 u_cpu.rf_ram.memory\[117\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09026__A2 _03962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09139_ _03134_ _04040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_68_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08785__A1 _03761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07588__A2 _03037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12150_ _00833_ net397 u_cpu.rf_ram.memory\[116\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10592__A1 _05053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11101_ u_cpu.cpu.genblk3.csr.mcause3_0\[3\] _05428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_78_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12081_ _00764_ net410 u_cpu.rf_ram.memory\[120\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06891__S0 _01651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[2\]_D net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08537__A1 _03588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11032_ _05379_ _05384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06012__A2 _01626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10895__A2 _05290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07760__A2 _03158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10647__A2 _05132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11934_ _00630_ net333 u_cpu.rf_ram.memory\[22\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11468__CLK net302 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11865_ _00561_ net519 u_cpu.rf_ram.memory\[136\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10816_ _05204_ _05245_ _05248_ _01176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08275__I _03490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11796_ _00492_ net374 u_cpu.rf_ram.memory\[73\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06079__A2 _01694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07276__A1 _02773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10747_ _04813_ _05204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10678_ u_cpu.rf_ram.memory\[102\]\[7\] _05150_ _05161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09017__A2 _03959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12417_ _01096_ net357 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05848__B _01455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout118_I net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07579__A2 _03036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12348_ _01027_ net117 u_cpu.rf_ram.memory\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10583__A1 _05044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10045__I _04737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12279_ _00962_ net525 u_arbiter.i_wb_cpu_dbus_adr\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08528__A1 _03602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout487_I net489 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07200__A1 _02726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06840_ _02078_ _02449_ _02450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06634__S0 _01779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10886__A2 _05293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06398__C _01900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06771_ u_cpu.rf_ram.memory\[44\]\[6\] u_cpu.rf_ram.memory\[45\]\[6\] u_cpu.rf_ram.memory\[46\]\[6\]
+ u_cpu.rf_ram.memory\[47\]\[6\] _01721_ _01624_ _02382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_114_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05762__A1 _01412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08510_ _03640_ _00477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05722_ u_cpu.cpu.csr_d_sel _01371_ _01372_ _01373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09490_ u_cpu.rf_ram.memory\[116\]\[5\] _04262_ _04266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08700__A1 u_cpu.rf_ram.memory\[137\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07503__A2 _02985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08441_ u_cpu.rf_ram.memory\[142\]\[3\] _03596_ _03599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08372_ _03494_ _03549_ _03554_ _00425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_17_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07323_ _02861_ u_cpu.rf_ram.memory\[1\]\[3\] _02852_ _02862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07267__A1 u_cpu.rf_ram.memory\[18\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05817__A2 _01461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07254_ _02768_ _02807_ _02814_ _00047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10810__A2 _05243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09008__A2 _03950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07019__A1 u_cpu.cpu.immdec.imm31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06205_ u_cpu.rf_ram.memory\[140\]\[0\] u_cpu.rf_ram.memory\[141\]\[0\] u_cpu.rf_ram.memory\[142\]\[0\]
+ u_cpu.rf_ram.memory\[143\]\[0\] _01820_ _01821_ _01822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07185_ _02762_ _02763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10949__I0 _04194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07529__I _03006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08767__A1 _03763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06136_ _01706_ _01753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10574__A1 _01443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06067_ _01683_ _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08519__A1 _03593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09744__I _04425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout401 net402 net401 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_47_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07990__A2 _03310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout412 net413 net412 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_132_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout423 net424 net423 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_113_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout434 net435 net434 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout445 net446 net445 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout456 net457 net456 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_09826_ u_arbiter.i_wb_cpu_rdt\[20\] u_arbiter.i_wb_cpu_rdt\[4\] _01442_ _04543_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06625__S0 _02029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout467 net473 net467 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout478 net484 net478 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_74_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout489 net493 net489 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09757_ _04464_ _04481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06969_ _01394_ _02576_ _02577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08708_ _02803_ _03380_ _03765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09688_ _01437_ _04413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08639_ _03720_ _00526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06553__I0 u_cpu.rf_ram.memory\[136\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11650_ _00354_ net216 u_cpu.rf_ram.memory\[60\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout30 net31 net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__11760__CLK net479 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09247__A2 _04109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout41 net42 net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_54_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10601_ _05113_ _01096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07258__A1 _02778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout52 net55 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_54_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11581_ _00285_ net339 u_cpu.rf_ram.memory\[68\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11054__A2 _05392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout63 net65 net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout74 net75 net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout85 net89 net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_126_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10532_ _05071_ _05072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout96 net97 net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__10801__A2 _05236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12116__CLK net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10463_ _04494_ _05021_ _05022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12202_ _00885_ net360 u_cpu.cpu.decode.opcode\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10394_ _04976_ _01026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10565__A1 u_cpu.rf_ram.memory\[96\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12133_ _00816_ net436 u_cpu.rf_ram.memory\[122\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12266__CLK net521 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07981__A2 _03303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12064_ _00747_ net289 u_cpu.rf_ram.memory\[35\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11015_ u_cpu.rf_ram.memory\[86\]\[3\] _05372_ _05374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10868__A2 _05270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08930__A1 u_cpu.rf_ram.memory\[128\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07733__A2 _03142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05744__A1 u_cpu.cpu.decode.op21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07902__I _03253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09486__A2 _04262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07497__A1 _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11917_ _00613_ net458 u_cpu.rf_ram.memory\[130\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11293__A2 _05548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07123__B _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11848_ _00544_ net509 u_cpu.rf_ram.memory\[137\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09238__A2 _04106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11045__A2 _02877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout235_I net240 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11779_ _00475_ net153 u_cpu.rf_ram.memory\[13\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06962__B _02564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09829__I _04450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08997__A1 u_cpu.rf_ram.memory\[125\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout402_I net414 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12609__CLK net380 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06224__A2 _01839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07421__A1 _02910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08990_ u_cpu.rf_ram.memory\[126\]\[7\] _03933_ _03944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07972__A2 _03300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07941_ _03264_ _03274_ _03281_ _00267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11746__D _00003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09174__A1 u_cpu.rf_ram.memory\[90\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07872_ _03193_ _03229_ _03236_ _00243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08221__I0 _02867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06527__A3 _02140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08921__A1 u_cpu.rf_ram.memory\[128\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07724__A2 _02891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09611_ _04356_ _04357_ _00862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06823_ u_cpu.rf_ram.memory\[128\]\[6\] u_cpu.rf_ram.memory\[129\]\[6\] u_cpu.rf_ram.memory\[130\]\[6\]
+ u_cpu.rf_ram.memory\[131\]\[6\] _01614_ _01616_ _02434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__11108__I0 u_cpu.cpu.genblk3.csr.mstatus_mie vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06083__S1 _01699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09542_ _03125_ net36 u_arbiter.i_wb_cpu_dbus_dat\[2\] _04286_ _04305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_110_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06754_ _02081_ _02364_ _01970_ _02365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11783__CLK net352 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06856__C _01427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09473_ _03918_ _04255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_36_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06685_ u_cpu.rf_ram.memory\[36\]\[5\] u_cpu.rf_ram.memory\[37\]\[5\] u_cpu.rf_ram.memory\[38\]\[5\]
+ u_cpu.rf_ram.memory\[39\]\[5\] _01716_ _02109_ _02297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_64_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08424_ _03586_ _00445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_u_scanchain_local.scan_flop\[26\]_D u_arbiter.i_wb_cpu_rdt\[23\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09229__A2 _04097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11036__A2 _05380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12139__CLK net398 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08355_ u_cpu.rf_ram.memory\[53\]\[4\] _03541_ _03544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07306_ _02725_ _02847_ _02848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08286_ _03498_ _03487_ _03499_ _00394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10795__A1 _05204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07237_ _02716_ _02782_ _02803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_20_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06302__I3 u_cpu.rf_ram.memory\[91\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06463__A2 _02070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07660__A1 _03071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09675__S _01438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12289__CLK net500 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09937__B1 _04502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06163__I _01632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07168_ _02726_ _02748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10547__A1 u_cpu.rf_ram.memory\[95\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06119_ _01685_ _01736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__07412__A1 _02897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07099_ _02675_ _02627_ _02686_ _02688_ _02689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_79_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout220 net221 net220 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout231 net268 net231 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_47_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout242 net246 net242 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout253 net254 net253 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout264 net265 net264 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout275 net281 net275 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout286 net288 net286 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__08912__A1 u_cpu.rf_ram.memory\[22\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09809_ _04526_ _04479_ _04528_ _04529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_8_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout297 net298 net297 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_21_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08818__I _03834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09468__A2 _04245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09712__I0 u_arbiter.i_wb_cpu_rdt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11702_ _00406_ net416 u_cpu.rf_ram.memory\[55\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_u_scanchain_local.scan_flop\[17\]_D u_arbiter.i_wb_cpu_rdt\[14\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12682_ _01360_ net100 u_cpu.rf_ram.memory\[23\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11633_ _00337_ net175 u_cpu.rf_ram.memory\[62\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08553__I _03484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11506__CLK net326 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11564_ _00268_ net343 u_cpu.rf_ram.memory\[75\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10786__A1 _05215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09640__A2 _04326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10515_ _05039_ _05060_ _05062_ _01061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07651__A1 _02723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11495_ _00199_ net99 u_cpu.rf_ram.memory\[17\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10446_ u_cpu.cpu.immdec.imm11_7\[1\] _04636_ _05005_ _05007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_137_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10377_ u_cpu.rf_ram.memory\[109\]\[3\] _04965_ _04967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12116_ _00799_ net116 u_cpu.rf_ram.memory\[11\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09156__A1 _03977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12047_ _00730_ net500 u_cpu.cpu.bufreg2.i_cnt_done vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout185_I net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10710__A1 _05137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09459__A2 _04245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07632__I _03074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout352_I net354 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11266__A2 _05527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11154__I _05464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08131__A2 _03394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06470_ _01573_ _02084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06142__A1 _01423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10993__I _02762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11018__A2 _05368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07890__A1 _03191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08140_ _03059_ _03405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09631__A2 _04285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08071_ _03347_ _03356_ _03363_ _00315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07642__A1 _03081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07079__I _02556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07022_ u_cpu.cpu.state.o_cnt\[2\] u_cpu.cpu.mem_bytecnt\[0\] _02628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__10529__A1 u_cpu.rf_ram.memory\[94\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08198__A2 _03439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12581__CLK net168 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout98_I net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07807__I _03080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07945__A2 _03275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08973_ _03933_ _03934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09147__A1 _02731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07924_ _03086_ _03270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[31\]_SE net547 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09698__A2 u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07855_ _03197_ _03217_ _03225_ _00237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10701__A1 _03165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06867__B _02476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06806_ _02150_ _02416_ _02153_ _02417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_44_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07786_ _03059_ _03179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_84_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09525_ _03132_ _04290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06771__I3 u_cpu.rf_ram.memory\[47\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06737_ u_cpu.rf_ram.memory\[132\]\[5\] u_cpu.rf_ram.memory\[133\]\[5\] u_cpu.rf_ram.memory\[134\]\[5\]
+ u_cpu.rf_ram.memory\[135\]\[5\] _02061_ _02174_ _02349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11529__CLK net488 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06133__A1 _01746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09456_ _04242_ _04239_ _04243_ _00821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06668_ _01590_ _02279_ _02280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09870__A2 _04526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08407_ _03576_ u_cpu.rf_ram.memory\[9\]\[7\] _03561_ _03577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06523__I3 u_cpu.rf_ram.memory\[119\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11009__A2 _05368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06684__A2 _02295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09607__C1 _04327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10609__S _05117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09387_ _04200_ u_cpu.rf_ram.memory\[8\]\[7\] _04185_ _04201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06599_ u_cpu.rf_ram.memory\[32\]\[4\] u_cpu.rf_ram.memory\[33\]\[4\] u_cpu.rf_ram.memory\[34\]\[4\]
+ u_cpu.rf_ram.memory\[35\]\[4\] _01705_ _01994_ _02212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_51_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05997__I _01613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08338_ _03504_ _03526_ _03533_ _00412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09622__A2 _04293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10768__A1 _05217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11679__CLK net314 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08269_ _03380_ _03166_ _03486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10300_ u_cpu.cpu.ctrl.o_ibus_adr\[6\] _04915_ _04917_ u_cpu.cpu.ctrl.o_ibus_adr\[7\]
+ _04919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_119_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11280_ u_cpu.rf_ram.memory\[89\]\[3\] _05539_ _05541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10231_ u_arbiter.i_wb_cpu_dbus_adr\[24\] u_arbiter.i_wb_cpu_dbus_adr\[23\] _04873_
+ _04875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_49_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08189__A2 _03310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06819__S0 _01831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07936__A2 _03278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10162_ _04835_ _04836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_120_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09138__A1 _02563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10093_ _04447_ _04774_ _04776_ _04779_ _04511_ _04780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__09932__I u_cpu.cpu.immdec.imm24_20\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12304__CLK net500 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06372__A1 _01876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10995_ _05359_ _05349_ _05360_ _01243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09310__A1 _04150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06068__I _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12454__CLK net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09861__A2 _04563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07872__A1 _03193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12665_ _01344_ net88 u_cpu.rf_ram.memory\[100\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08283__I _02756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11616_ _00320_ net101 u_cpu.rf_ram.memory\[29\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10759__A1 _05211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12596_ _01275_ net274 u_cpu.rf_ram.memory\[88\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10318__I _04905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06427__A2 _02041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07624__A1 u_cpu.rf_ram.memory\[47\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07120__C _02705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11547_ _00251_ net258 u_cpu.rf_ram.memory\[74\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11478_ _00182_ net121 u_cpu.rf_ram.memory\[4\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout100_I net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10429_ _04814_ _04993_ _04996_ _01041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[54\]_SE net561 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07627__I _03070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06286__S1 _01737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10931__A1 u_cpu.rf_ram.memory\[59\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11149__I _02777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05970_ _01417_ _01587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08352__A2 _03537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07640_ _03080_ _03081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06363__A1 _01649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07362__I _02739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07571_ _02875_ _02936_ _03033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__11239__A2 _05511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06753__I3 u_cpu.rf_ram.memory\[19\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09310_ _04150_ _04142_ _04151_ _00767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06522_ _01704_ _02136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_74_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09852__A2 _04567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10998__A1 _05361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06453_ _01570_ _02066_ _02067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09241_ _04061_ _04105_ _04108_ _00741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07863__A1 _03179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09172_ _04056_ _04058_ _04060_ _00719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout13_I net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06384_ _01862_ _01985_ _01998_ _01999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_119_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09604__A2 _04352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08123_ u_cpu.rf_ram.memory\[62\]\[0\] _03395_ _03396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10228__I _02690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06269__I2 u_cpu.rf_ram.memory\[34\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08054_ _03351_ _03338_ _03352_ _00309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07091__A2 _02680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07005_ _02610_ _02611_ _02612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_31_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08415__I0 _03566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05929__A1 _01524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06277__S1 _01892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10922__A1 u_cpu.rf_ram.memory\[59\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12327__CLK net525 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08591__A2 _03691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08956_ _03894_ _03922_ _03924_ _00639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07907_ _03257_ _03254_ _03258_ _00256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10898__I _02730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08887_ _03876_ _00618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08343__A2 _03425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07838_ _03033_ _03202_ _03215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11351__CLK net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07769_ u_cpu.rf_ram.memory\[40\]\[0\] _03169_ _03170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09508_ u_cpu.rf_ram.memory\[33\]\[4\] _04274_ _04277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_77_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10780_ _05209_ _05220_ _05226_ _01162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10989__A1 _05354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06657__A2 _02268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09439_ _04150_ _04226_ _04232_ _00815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12450_ _01129_ net87 u_cpu.rf_ram.memory\[103\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11401_ _00105_ net294 u_cpu.rf_ram.memory\[42\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10138__I _04809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07606__A1 _02994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12381_ _01060_ net76 u_cpu.rf_ram.memory\[97\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11332_ _00036_ net59 u_cpu.rf_ram.memory\[21\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07082__A2 u_cpu.cpu.state.o_cnt_r\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11263_ _02906_ _05523_ _05530_ _01341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10214_ _04865_ _00957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08031__A1 _02804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11194_ _05488_ _05490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10913__A1 u_cpu.rf_ram.memory\[84\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10145_ _02761_ _04823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10076_ _04420_ _04455_ _04604_ _04764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_48_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09531__A1 u_arbiter.i_wb_cpu_rdt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08334__A2 _03525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08278__I _02750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11844__CLK net421 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08098__A1 _03353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10978_ _02920_ _05243_ _05348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06648__A2 _02260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout148_I net156 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12648_ _01327_ net142 u_cpu.rf_ram.memory\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11994__CLK net259 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09598__A1 u_arbiter.i_wb_cpu_rdt\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout315_I net323 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12579_ _01258_ net166 u_cpu.rf_ram.memory\[111\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10904__A1 u_cpu.rf_ram.memory\[84\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08573__A2 _03674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08810_ _03828_ _03817_ _03829_ _00588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09790_ _04416_ _04510_ _04447_ _04423_ _04511_ _04512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_100_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11374__CLK net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10380__A2 _04961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05926__A4 _01535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08741_ _03757_ _03778_ _03785_ _00563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05953_ _01569_ _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_94_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05884_ _01473_ _01514_ _01515_ u_arbiter.o_wb_cpu_adr\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08672_ u_cpu.rf_ram.memory\[39\]\[4\] _03738_ _03741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07623_ _03067_ _03068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_81_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08916__I _02738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07554_ u_cpu.rf_ram.memory\[41\]\[0\] _03023_ _03024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09825__A2 _04396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06505_ _02117_ _02118_ _02119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06639__A2 _02251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07836__A1 u_cpu.rf_ram.memory\[129\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07485_ _02904_ _02969_ _02975_ _00117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08884__I0 _03566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09224_ _04063_ _04093_ _04098_ _00734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06436_ _02042_ _02044_ _02046_ _02049_ _02050_ _02051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_21_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08636__I0 _03574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09155_ u_cpu.rf_ram.memory\[91\]\[2\] _04049_ _04050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06367_ _01666_ _01981_ _01982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06880__B _01679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08106_ _03340_ _03382_ _03385_ _00328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07064__A2 _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06298_ _01423_ _01901_ _01913_ _01914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_09086_ u_cpu.rf_ram.memory\[37\]\[1\] _04004_ _04006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08037_ u_cpu.rf_ram.memory\[65\]\[1\] _03338_ _03341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06811__A2 _02421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11148__A1 _05460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11717__CLK net417 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06171__I _01575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08564__A2 _03674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09988_ _04684_ _04685_ _00911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10371__A2 _04961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08939_ _03910_ _03896_ _03911_ _00635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11867__CLK net519 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09513__A1 _04253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08316__A2 _03513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11950_ _00646_ net451 u_cpu.rf_ram.memory\[127\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10123__A2 u_cpu.cpu.genblk3.csr.mstatus_mie vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11320__A1 _03119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10901_ _05301_ _05303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06878__A2 _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11881_ _00577_ net518 u_cpu.rf_ram.memory\[134\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10832_ _05256_ _05258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09816__A2 _04457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07827__A1 _03188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10763_ _04829_ _05215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_41_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11252__I _05522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12502_ _01181_ net39 u_cpu.rf_ram.memory\[107\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10694_ _05142_ _05164_ _05171_ _01131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12433_ _01112_ net160 u_cpu.rf_ram.memory\[101\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12364_ _01043_ net210 u_cpu.rf_ram.memory\[93\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11315_ _02648_ u_cpu.rf_ram.rdata\[7\] u_cpu.rf_ram_if.rtrig0 _05561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_107_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[39\] u_scanchain_local.module_data_in\[38\] net552 u_arbiter.o_wb_cpu_adr\[1\]
+ net20 u_scanchain_local.module_data_in\[39\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__11139__A1 _05454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12295_ _00977_ net93 u_cpu.rf_ram.memory\[30\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11397__CLK net299 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06081__I _01650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12642__CLK net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11246_ u_cpu.rf_ram.memory\[98\]\[6\] _05515_ _05520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06405__I2 u_cpu.rf_ram.memory\[114\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11177_ u_cpu.rf_ram.memory\[25\]\[1\] _05478_ _05480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07905__I _03067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10128_ _04809_ _04810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09504__A1 u_cpu.rf_ram.memory\[33\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08307__A2 _03513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10059_ _04509_ _04548_ _04748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07126__B u_cpu.rf_ram_if.genblk1.wtrig0_r vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10114__A2 _02625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout265_I net266 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07640__I _03080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07818__A1 _02804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout432_I net433 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06177__S0 _01792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07270_ _02758_ _02818_ _02824_ _00053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07294__A2 _02837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06097__A3 _01646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06221_ _01564_ _01714_ _01837_ _00000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__12172__CLK net386 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[31\]_CLK net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06152_ u_cpu.rf_ram.memory\[88\]\[0\] u_cpu.rf_ram.memory\[89\]\[0\] u_cpu.rf_ram.memory\[90\]\[0\]
+ u_cpu.rf_ram.memory\[91\]\[0\] _01767_ _01768_ _01769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_121_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11749__D _00006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09991__A1 _04497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06083_ u_cpu.rf_ram.memory\[36\]\[0\] u_cpu.rf_ram.memory\[37\]\[0\] u_cpu.rf_ram.memory\[38\]\[0\]
+ u_cpu.rf_ram.memory\[39\]\[0\] _01698_ _01699_ _01700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08794__A2 _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09911_ _04610_ _04616_ _04617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_u_scanchain_local.scan_flop\[46\]_CLK net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08546__A2 _03655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09842_ _04498_ _04558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout80_I net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09516__B _04031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06101__S0 _01716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09773_ _04484_ _04485_ _04488_ _04495_ _04496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_80_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06985_ _01385_ u_cpu.cpu.state.init_done _01386_ _01376_ _02592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08724_ u_cpu.rf_ram.memory\[49\]\[6\] _03770_ _03775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05936_ u_arbiter.i_wb_cpu_dbus_adr\[29\] _01493_ _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10105__A2 _04788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11302__A1 u_cpu.rf_ram.memory\[23\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08655_ _03680_ _03723_ _03730_ _00532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05867_ u_cpu.cpu.ctrl.o_ibus_adr\[14\] _01502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06875__B _01663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07606_ _02994_ _03048_ _03055_ _00158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08586_ u_cpu.rf_ram.memory\[70\]\[1\] _03688_ _03690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05798_ _01443_ _01444_ _01445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07550__I _03019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07809__A1 _03195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07537_ _02989_ _03007_ _03012_ _00132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_41_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07468_ _02913_ _02955_ _02963_ _00112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06332__I1 u_cpu.rf_ram.memory\[129\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09207_ _02557_ _04086_ _04087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_52_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06419_ u_cpu.rf_ram.memory\[80\]\[2\] u_cpu.rf_ram.memory\[81\]\[2\] u_cpu.rf_ram.memory\[82\]\[2\]
+ u_cpu.rf_ram.memory\[83\]\[2\] _01773_ _02033_ _02034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_52_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10617__S _05117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06883__I2 u_cpu.rf_ram.memory\[118\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07399_ _02916_ _02894_ _02917_ _00089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07037__A2 _02640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09138_ _02563_ _04038_ _04039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10041__A1 _04732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10041__B2 _04467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08785__A2 _03803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09069_ u_cpu.rf_ram.memory\[38\]\[2\] _03995_ _03996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06796__A1 _01691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06115__B _01731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11100_ _05418_ _05426_ _05427_ _01281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_12080_ _00763_ net312 u_cpu.rf_ram.memory\[117\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06891__S1 _01653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08537__A2 _03655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11031_ _05352_ _05380_ _05383_ _01256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_46_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06643__S1 _01942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12045__CLK net495 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07348__I0 _02855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09940__I _04489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11933_ _00629_ net419 u_cpu.rf_ram.memory\[22\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11864_ _00560_ net517 u_cpu.rf_ram.memory\[136\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12195__CLK net398 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10815_ u_cpu.rf_ram.memory\[107\]\[1\] _05246_ _05248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11795_ _00491_ net373 u_cpu.rf_ram.memory\[73\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06076__I _01659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07276__A2 _02819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10746_ _05199_ _05201_ _05203_ _01151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_41_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10280__A1 _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10677_ _05146_ _05152_ _05160_ _01125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10407__I0 _04184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12416_ _01095_ net357 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07028__A2 u_cpu.cpu.decode.opcode\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08291__I _02766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10032__A1 _04721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08776__A2 _03806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12347_ _01026_ net116 u_cpu.rf_ram.memory\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12278_ _00961_ net532 u_arbiter.i_wb_cpu_dbus_adr\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08528__A2 _03644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11229_ _05509_ _01328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07635__I _02762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07200__A2 u_cpu.rf_ram_if.wdata1_r\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06634__S1 _01930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout382_I net393 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06770_ _01772_ _02380_ _02381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07339__I0 _02873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05762__A2 _01377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10099__A1 _04548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05721_ u_cpu.cpu.bne_or_bge _01372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_82_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10996__I _02767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11412__CLK net226 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06695__B _01587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12538__CLK net279 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08440_ _03497_ _03598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08700__A2 _03753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08371_ u_cpu.rf_ram.memory\[52\]\[2\] _03553_ _03554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10010__B _04704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07322_ _02860_ _02861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11562__CLK net259 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08464__A1 _03595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07267__A2 _02822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12688__CLK net234 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10271__A1 _04821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07253_ u_cpu.rf_ram.memory\[81\]\[5\] _02810_ _02814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06570__S0 _01959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09297__I _04141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06204_ _01815_ _01821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_121_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07184_ _02761_ _02762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10023__A1 _04715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09964__A1 _04585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06135_ _01704_ _01752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08767__A2 _03791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06778__A1 _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06066_ _01568_ _01683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08519__A2 _03643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout402 net414 net402 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_28_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout413 net414 net413 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12068__CLK net282 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout424 net434 net424 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__10326__A2 _04929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout435 net476 net435 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_58_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout446 net447 net446 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_115_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09825_ _01409_ _04396_ _04542_ _00891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout457 net459 net457 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_63_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout468 net469 net468 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_101_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06625__S1 _01742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout479 net483 net479 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_58_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09756_ _04468_ _04469_ _04479_ _04480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06968_ _01411_ _02555_ _02558_ _02560_ _02575_ _02576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XANTENNA__06950__A1 _02556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08707_ _03763_ _03748_ _03764_ _00550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05919_ u_arbiter.i_wb_cpu_dbus_adr\[25\] _01539_ _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09687_ _04409_ _04411_ _04412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06899_ _01778_ _02508_ _01782_ _02509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08638_ _03576_ u_cpu.rf_ram.memory\[14\]\[7\] _03711_ _03720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06553__I1 u_cpu.rf_ram.memory\[137\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11905__CLK net471 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08569_ _03500_ _03678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_126_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout20 net25 net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout31 net32 net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_70_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10600_ u_arbiter.i_wb_cpu_rdt\[17\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\]
+ _05111_ _05113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xfanout42 net43 net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__07258__A2 _02807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout53 net55 net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__08455__A1 _02966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11580_ _00284_ net340 u_cpu.rf_ram.memory\[68\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout64 net65 net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_126_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout75 net78 net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_50_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout86 net89 net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_50_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10531_ _04091_ _03062_ _05071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout97 net100 net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_52_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06561__S0 _02061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08207__A1 u_cpu.rf_ram.memory\[19\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10462_ _04444_ _05018_ _05020_ _04747_ _05021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_13_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10014__A1 _04477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12201_ _00884_ net384 u_cpu.cpu.decode.opcode\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09955__A1 _04585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08758__A2 _03794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06608__I2 u_cpu.rf_ram.memory\[102\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10393_ _04190_ u_cpu.rf_ram.memory\[3\]\[2\] _04973_ _04976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10565__A2 _05088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12132_ _00815_ net436 u_cpu.rf_ram.memory\[122\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12063_ _00746_ net307 u_cpu.rf_ram.memory\[35\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11014_ _05354_ _05368_ _05373_ _01249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07194__A1 _02748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11435__CLK net334 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08930__A2 _03904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06941__A1 _02549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11916_ _00612_ net454 u_cpu.rf_ram.memory\[130\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11585__CLK net248 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08694__A1 u_cpu.rf_ram.memory\[137\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07497__A2 _02982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07190__I _02766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11847_ _00543_ net508 u_cpu.rf_ram.memory\[137\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10628__I0 u_arbiter.i_wb_cpu_rdt\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07249__A2 _02810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11778_ _00474_ net152 u_cpu.rf_ram.memory\[13\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10253__A1 _02690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08997__A2 _03947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout130_I net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10729_ u_cpu.rf_ram.memory\[99\]\[2\] _05192_ _05193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout228_I net229 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09946__A1 u_cpu.cpu.immdec.imm24_20\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06304__S0 _01773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12210__CLK net352 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07421__A2 _02926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07940_ u_cpu.rf_ram.memory\[75\]\[4\] _03278_ _03281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07365__I _02890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09174__A2 _04059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07871_ u_cpu.rf_ram.memory\[77\]\[4\] _03233_ _03236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09610_ u_arbiter.i_wb_cpu_rdt\[18\] _04347_ _04344_ u_arbiter.i_wb_cpu_dbus_dat\[18\]
+ _04357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_68_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08921__A2 _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06822_ _01830_ _02432_ _01628_ _02433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06932__A1 u_cpu.cpu.bufreg2.i_cnt_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11928__CLK net333 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09541_ u_arbiter.i_wb_cpu_dbus_dat\[3\] _04286_ _04304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_23_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06753_ u_cpu.rf_ram.memory\[16\]\[6\] u_cpu.rf_ram.memory\[17\]\[6\] u_cpu.rf_ram.memory\[18\]\[6\]
+ u_cpu.rf_ram.memory\[19\]\[6\] _01598_ _01968_ _02364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_77_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09472_ _04253_ _04240_ _04254_ _00826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout43_I net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07488__A2 _02973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08196__I _03438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08685__A1 _03745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06684_ _01988_ _02295_ _02107_ _02296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_58_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08423_ _03574_ u_cpu.rf_ram.memory\[15\]\[6\] _03578_ _03586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06791__S0 _01674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08354_ _03498_ _03537_ _03543_ _00418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08924__I _03899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07305_ u_cpu.cpu.immdec.imm11_7\[3\] _02724_ _02847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08988__A2 _03938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08285_ u_cpu.rf_ram.memory\[56\]\[3\] _03495_ _03499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10795__A2 _05232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07236_ _02778_ _02793_ _02802_ _00041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07660__A2 _03090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09937__A1 _04549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07167_ _02733_ _02746_ _02747_ _00027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10547__A2 _05076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06118_ _01648_ _01735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_65_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07412__A2 _02925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07098_ u_cpu.cpu.bufreg.c_r _02687_ _02688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_79_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06471__I0 u_cpu.rf_ram.memory\[28\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12703__CLK net235 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06049_ _01665_ _01666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout210 net211 net210 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_82_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout221 net223 net221 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout232 net235 net232 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__09165__A2 _04044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout243 net244 net243 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_47_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout254 net255 net254 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout265 net266 net265 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__07176__A1 _02748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout276 net280 net276 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_09808_ _04527_ _04528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout287 net288 net287 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__08912__A2 _03886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10630__S _03116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout298 net305 net298 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09739_ _04404_ u_arbiter.i_wb_cpu_ibus_adr\[1\] _04463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07479__A2 _02970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08676__A1 u_cpu.rf_ram.memory\[39\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11701_ _00405_ net415 u_cpu.rf_ram.memory\[55\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12681_ _01359_ net97 u_cpu.rf_ram.memory\[23\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06782__S0 _02005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11632_ _00336_ net175 u_cpu.rf_ram.memory\[62\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08428__A1 _02920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09625__B1 _04359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11563_ _00267_ net341 u_cpu.rf_ram.memory\[75\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06534__S0 _01773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10786__A2 _05221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10514_ u_cpu.rf_ram.memory\[94\]\[0\] _05061_ _05062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12233__CLK net359 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11494_ _00198_ net98 u_cpu.rf_ram.memory\[16\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07651__A2 _03005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09928__A1 _04629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10445_ _05005_ _05006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08600__A1 _03684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10376_ _04817_ _04961_ _04966_ _01018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_48_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[21\] u_arbiter.i_wb_cpu_rdt\[18\] net541 u_arbiter.i_wb_cpu_dbus_dat\[15\]
+ net9 u_arbiter.i_wb_cpu_rdt\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
X_12115_ _00798_ net116 u_cpu.rf_ram.memory\[11\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06303__B _01770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07185__I _02762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12046_ _00729_ net495 u_cpu.cpu.ctrl.i_jump vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07118__C _02605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07167__A1 _02733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06914__A1 _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10710__A2 _05176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout345_I net356 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06142__A2 _01734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06773__S0 _01716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07890__A2 _03241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout512_I net514 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09092__A1 _03980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10777__A2 _05224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08070_ u_cpu.rf_ram.memory\[64\]\[4\] _03360_ _03363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09919__A1 _04620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07021_ _02569_ _02625_ _02626_ _02627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11600__CLK net244 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10529__A2 _05059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08972_ _02920_ _03181_ _03933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11750__CLK net254 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07923_ _03268_ _03255_ _03269_ _00261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09147__A2 _03034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07854_ u_cpu.rf_ram.memory\[139\]\[6\] _03220_ _03225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08919__I _03895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06905__A1 _01565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10701__A2 _05162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06805_ u_cpu.rf_ram.memory\[84\]\[6\] u_cpu.rf_ram.memory\[85\]\[6\] u_cpu.rf_ram.memory\[86\]\[6\]
+ u_cpu.rf_ram.memory\[87\]\[6\] _01752_ _02151_ _02416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_72_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12106__CLK net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07785_ _03087_ _03169_ _03178_ _00214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09524_ _03124_ _04289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08658__A1 u_cpu.rf_ram.memory\[138\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06736_ _01947_ _02347_ _02348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_77_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10465__A1 _04518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09455_ u_cpu.rf_ram.memory\[115\]\[1\] _04240_ _04243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06667_ u_cpu.rf_ram.memory\[28\]\[5\] u_cpu.rf_ram.memory\[29\]\[5\] u_cpu.rf_ram.memory\[30\]\[5\]
+ u_cpu.rf_ram.memory\[31\]\[5\] _02084_ _01577_ _02279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06133__A2 _01749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08406_ _02872_ _03576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_40_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09607__B1 _04321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09386_ _02872_ _04200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_75_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12256__CLK net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06598_ _01882_ _02210_ _02211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05892__A1 _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08337_ u_cpu.rf_ram.memory\[54\]\[5\] _03529_ _03533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06174__I _01777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08830__A1 _03826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08268_ _03484_ _03485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07633__A2 _03072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06692__I0 u_cpu.rf_ram.memory\[108\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07219_ _02791_ _02793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08199_ u_cpu.rf_ram.memory\[19\]\[3\] _03443_ _03445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10230_ _04874_ _00964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06819__S1 _01832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10424__I _04992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10161_ _03367_ _03062_ _04835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10092_ _04692_ _04751_ _04778_ _04575_ _04779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_48_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06777__C _01733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08649__A1 _03673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10994_ u_cpu.rf_ram.memory\[110\]\[4\] _05355_ _05360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10456__A1 _04680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09310__A2 _04142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10456__B2 _04482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06755__S0 _02084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12664_ _01343_ net86 u_cpu.rf_ram.memory\[100\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07872__A2 _03229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11615_ _00319_ net101 u_cpu.rf_ram.memory\[29\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09074__A1 _03982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11623__CLK net185 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[69\] u_scanchain_local.module_data_in\[68\] net559 u_arbiter.o_wb_cpu_adr\[31\]
+ net27 u_scanchain_local.module_data_in\[69\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
X_12595_ _01274_ net274 u_cpu.rf_ram.memory\[88\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10759__A2 _05201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11546_ _00250_ net258 u_cpu.rf_ram.memory\[74\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08821__A1 _03813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11477_ _00181_ net67 u_cpu.rf_ram.memory\[4\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07908__I _03070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11773__CLK net514 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10428_ u_cpu.rf_ram.memory\[93\]\[1\] _04994_ _04996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11184__A2 _05481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10359_ _04952_ _02579_ _04953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10931__A2 _05318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12129__CLK net410 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout295_I net298 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12029_ _00712_ net313 u_cpu.rf_ram.memory\[91\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07643__I _02772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout462_I net467 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06363__A2 _01977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07560__A1 _02989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07570_ _03000_ _03023_ _03032_ _00145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12279__CLK net525 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10447__A1 _02535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06521_ _01746_ _02134_ _02135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10447__B2 _04732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06115__A2 _01730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06746__S0 _01959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09240_ u_cpu.rf_ram.memory\[35\]\[1\] _04106_ _04108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06452_ u_cpu.rf_ram.memory\[8\]\[3\] u_cpu.rf_ram.memory\[9\]\[3\] u_cpu.rf_ram.memory\[10\]\[3\]
+ u_cpu.rf_ram.memory\[11\]\[3\] _01574_ _01838_ _02066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07863__A2 _03229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09171_ u_cpu.rf_ram.memory\[90\]\[0\] _04059_ _04060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09065__A1 _03969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06383_ _01987_ _01990_ _01992_ _01997_ _01711_ _01998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_08122_ _03393_ _03395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07615__A2 _02919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08053_ u_cpu.rf_ram.memory\[65\]\[6\] _03343_ _03352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07004_ u_arbiter.i_wb_cpu_ibus_adr\[0\] u_cpu.cpu.ctrl.pc_plus_4_cy_r _02611_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07379__A1 _02900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06426__I0 u_cpu.rf_ram.memory\[64\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11175__A2 _05478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08955_ u_cpu.rf_ram.memory\[127\]\[0\] _03923_ _03924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07906_ u_cpu.rf_ram.memory\[76\]\[1\] _03255_ _03258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08886_ _03568_ u_cpu.rf_ram.memory\[12\]\[3\] _03872_ _03876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_9_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07837_ _03199_ _03205_ _03214_ _00230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07551__A1 _03018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06169__I _01683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07768_ _03167_ _03169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09507_ _04247_ _04270_ _04276_ _00839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10438__A1 _04827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06719_ _02324_ _02326_ _02328_ _02330_ _01925_ _02331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_38_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11646__CLK net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07699_ _02569_ _02695_ _02598_ _03120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06737__S0 _02061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10989__A2 _05349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09438_ u_cpu.rf_ram.memory\[122\]\[3\] _04230_ _04232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07854__A2 _03220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05865__A1 _01489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09369_ _04188_ u_cpu.rf_ram.memory\[8\]\[1\] _04186_ _04189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_36_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11400_ _00104_ net293 u_cpu.rf_ram.memory\[42\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11796__CLK net374 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12380_ _01059_ net80 u_cpu.rf_ram.memory\[97\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07606__A2 _03048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11331_ _00035_ net68 u_cpu.rf_ram.memory\[21\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09359__A2 _04177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11262_ u_cpu.rf_ram.memory\[100\]\[4\] _05527_ _05530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11166__A2 _05469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10213_ u_arbiter.i_wb_cpu_dbus_adr\[16\] u_arbiter.i_wb_cpu_dbus_adr\[15\] _04861_
+ _04865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10154__I _04829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08031__A2 _02923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11193_ _05488_ _05489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_122_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10144_ _04821_ _04810_ _04822_ _00930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10075_ _04407_ _04709_ _04474_ _04763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08559__I _03490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09531__A2 _04293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10677__A1 _05146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10429__A1 _04814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10977_ _02739_ _05347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08098__A2 _03370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12571__CLK net200 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09834__A3 _04550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12647_ _01326_ net133 u_cpu.rf_ram.memory\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09047__A1 u_cpu.rf_ram.memory\[123\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06028__B _01644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09598__A2 _04326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12578_ _01257_ net172 u_cpu.rf_ram.memory\[111\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11529_ _00233_ net488 u_cpu.rf_ram.memory\[139\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout210_I net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout308_I net311 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06900__S0 _01762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06281__A1 _01725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11157__A2 _05466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08022__A2 _03328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11519__CLK net430 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10904__A2 _05303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10999__I _02772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07781__A1 _03081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08740_ u_cpu.rf_ram.memory\[136\]\[4\] _03782_ _03785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05952_ _01568_ _01569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_61_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10668__A1 u_cpu.rf_ram.memory\[102\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08671_ _03676_ _03734_ _03740_ _00538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05883_ u_arbiter.i_wb_cpu_dbus_adr\[17\] _01481_ _01515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11669__CLK net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06187__I2 u_cpu.rf_ram.memory\[78\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07622_ _02745_ _03067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07553_ _03021_ _03023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09286__A1 _04066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06504_ u_cpu.rf_ram.memory\[108\]\[3\] u_cpu.rf_ram.memory\[109\]\[3\] u_cpu.rf_ram.memory\[110\]\[3\]
+ u_cpu.rf_ram.memory\[111\]\[3\] _02001_ _01717_ _02118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_34_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07484_ u_cpu.rf_ram.memory\[45\]\[3\] _02973_ _02975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09223_ u_cpu.rf_ram.memory\[92\]\[2\] _04097_ _04098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06435_ _01606_ _02050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09038__A1 _03969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09154_ _04044_ _04049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08932__I _02756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06366_ u_cpu.rf_ram.memory\[60\]\[2\] u_cpu.rf_ram.memory\[61\]\[2\] u_cpu.rf_ram.memory\[62\]\[2\]
+ u_cpu.rf_ram.memory\[63\]\[2\] _01639_ _01668_ _01981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08105_ u_cpu.rf_ram.memory\[63\]\[1\] _03383_ _03385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09085_ _03969_ _04003_ _04005_ _00687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06297_ _01903_ _01907_ _01910_ _01912_ _01757_ _01913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__08261__A2 _03477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07548__I _02939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08036_ _03067_ _03340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_123_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09210__A1 _04034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08013__A2 _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10356__B1 _04909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09763__I _04472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12444__CLK net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09987_ u_cpu.cpu.immdec.imm30_25\[2\] _04672_ _04674_ u_cpu.cpu.immdec.imm30_25\[3\]
+ _04682_ _04558_ _04685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__07772__A1 _03068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10702__I _05175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08938_ u_cpu.rf_ram.memory\[128\]\[4\] _03904_ _03911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07283__I _02832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10659__A1 _05148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09513__A2 _04271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08869_ u_cpu.rf_ram.memory\[130\]\[4\] _03863_ _03866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07524__A1 _02716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10123__A3 u_cpu.cpu.genblk3.csr.i_mtip vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12594__CLK net279 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10900_ _05301_ _05302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_44_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11880_ _00576_ net456 u_cpu.rf_ram.memory\[134\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10831_ _05256_ _05257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11084__A1 _05365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10762_ _05213_ _05202_ _05214_ _01156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[44\]_SE net559 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12501_ _01180_ net39 u_cpu.rf_ram.memory\[107\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09029__A1 _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10149__I _02766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10693_ u_cpu.rf_ram.memory\[103\]\[4\] _05168_ _05171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12432_ _01111_ net88 u_cpu.rf_ram.memory\[101\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12363_ _01042_ net211 u_cpu.rf_ram.memory\[93\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08252__A2 _03474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11314_ _05560_ _01362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12294_ _00976_ net94 u_cpu.rf_ram.memory\[30\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11245_ _05458_ _05512_ _05519_ _01334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09201__A1 _02547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08004__A2 _03316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09673__I _04397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11176_ _05444_ _05477_ _05479_ _01305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07763__A1 _03087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11811__CLK net376 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10127_ _02890_ _02965_ _04809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10058_ _04692_ _04709_ _04474_ _04747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_23_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11311__A2 _05558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07921__I _03083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout160_I net164 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09268__A1 _04068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout258_I net259 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11075__A1 u_cpu.rf_ram.memory\[88\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06537__I _01632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07818__A2 _03202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06177__S1 _01793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05829__A1 u_cpu.cpu.ctrl.o_ibus_adr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12317__CLK net524 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout425_I net429 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08491__A2 _03625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06220_ _01811_ _01836_ _01837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06151_ _01675_ _01768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08243__A2 _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10050__A2 _04636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12467__CLK net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06082_ _01667_ _01699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10008__B _04703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09910_ _04567_ _04612_ _04615_ _04616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_99_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10338__B1 _04938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09583__I _04318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09841_ _01382_ _04396_ _04557_ _00892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10889__A1 _05278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06557__A2 _02170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07754__A1 u_cpu.rf_ram.memory\[17\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06101__S1 _01717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06801__I0 u_cpu.rf_ram.memory\[88\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09772_ _04484_ _04492_ _04494_ _04495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06984_ _01369_ _02591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_101_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout73_I net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08723_ _03759_ _03767_ _03774_ _00556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05935_ u_cpu.cpu.ctrl.o_ibus_adr\[29\] _01554_ _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_80_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08654_ u_cpu.rf_ram.memory\[138\]\[5\] _03726_ _03730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05866_ u_arbiter.i_wb_cpu_dbus_adr\[14\] _01453_ _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08927__I _02750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[67\]_SE net554 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07605_ u_cpu.rf_ram.memory\[48\]\[4\] _03052_ _03055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08585_ _03666_ _03687_ _03689_ _00503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09259__A1 _04056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05797_ u_cpu.cpu.ctrl.o_ibus_adr\[2\] _01444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_74_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07536_ u_cpu.rf_ram.memory\[51\]\[2\] _03011_ _03012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07467_ u_cpu.rf_ram.memory\[46\]\[6\] _02958_ _02963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09206_ _04083_ _04084_ _04085_ _02589_ _04086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06418_ _01652_ _02033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07398_ u_cpu.rf_ram.memory\[80\]\[7\] _02892_ _02917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06883__I3 u_cpu.rf_ram.memory\[119\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09137_ _04037_ _04038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06349_ _01955_ _01957_ _01961_ _01963_ _01607_ _01964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_33_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06182__I _01584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09068_ _03990_ _03995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08019_ _03259_ _03324_ _03329_ _00297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_78_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11030_ u_cpu.rf_ram.memory\[111\]\[1\] _05381_ _05383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11984__CLK net438 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11932_ _00628_ net333 u_cpu.rf_ram.memory\[22\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11863_ _00559_ net516 u_cpu.rf_ram.memory\[136\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10814_ _05199_ _05245_ _05247_ _01175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11794_ _00490_ net352 u_cpu.rf_ram.memory\[73\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10100__C _04459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10804__A1 _05213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10745_ u_cpu.rf_ram.memory\[79\]\[0\] _05202_ _05203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08473__A2 _03608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11364__CLK net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10280__A2 _02705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08572__I _03503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10676_ u_cpu.rf_ram.memory\[102\]\[6\] _05155_ _05160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12415_ _01094_ net82 u_cpu.rf_ram.memory\[28\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xu_scanchain_local.scan_flop\[51\] u_scanchain_local.module_data_in\[50\] net560 u_arbiter.o_wb_cpu_adr\[13\]
+ net29 u_scanchain_local.module_data_in\[51\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__09422__A1 _04154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10032__A2 _04489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12346_ _01025_ net117 u_cpu.rf_ram.memory\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06092__I _01662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09973__A2 _04672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07984__A1 _03266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06787__A2 _02397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12277_ _00960_ net533 u_arbiter.i_wb_cpu_dbus_adr\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09725__A2 u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.out_flop u_scanchain_local.module_data_in\[69\] net26 u_scanchain_local.data_out_i
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_11228_ _02872_ u_cpu.rf_ram.memory\[0\]\[7\] _05500_ _05509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10342__I _04905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11159_ _05464_ _05469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_fanout375_I net382 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09489__A1 _04249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05720_ u_cpu.cpu.decode.co_mem_word _01371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_23_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11296__A1 _02896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08161__A1 _03419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout542_I net546 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11173__I _05476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08370_ _03548_ _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07321_ u_cpu.rf_ram_if.wdata0_r\[3\] u_cpu.rf_ram_if.wdata1_r\[3\] _02844_ _02860_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_75_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08464__A2 _03609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09661__A1 _04247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08482__I _03620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10271__A2 _04894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07252_ _02763_ _02806_ _02813_ _00046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06203_ _01613_ _01820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06570__S1 _02071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07183_ _02735_ u_cpu.rf_ram_if.wdata0_r\[4\] _02760_ _02761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__09413__A1 _04145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11857__CLK net420 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06227__A1 _01580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06134_ _01609_ _01751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09964__A2 _04663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07975__A1 _03257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06065_ _01655_ _01664_ _01670_ _01680_ _01681_ _01682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__09716__A2 u_arbiter.i_wb_cpu_rdt\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout403 net407 net403 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_98_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout414 net435 net414 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout425 net429 net425 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_101_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout436 net442 net436 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_101_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09824_ _04516_ _04541_ _04542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout447 net448 net447 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout458 net459 net458 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout469 net472 net469 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06250__I1 u_cpu.rf_ram.memory\[49\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09755_ _04474_ _04478_ _04479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06967_ _02561_ _02545_ _02567_ u_cpu.cpu.genblk3.csr.mstatus_mie _02574_ _02575_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_104_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06950__A2 _02557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05918_ u_cpu.cpu.ctrl.o_ibus_adr\[25\] _01541_ _01542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08706_ u_cpu.rf_ram.memory\[137\]\[7\] _03746_ _03764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11287__A1 _02912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09686_ _04404_ u_arbiter.i_wb_cpu_rdt\[12\] _04410_ _04411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06898_ u_cpu.rf_ram.memory\[68\]\[7\] u_cpu.rf_ram.memory\[69\]\[7\] u_cpu.rf_ram.memory\[70\]\[7\]
+ u_cpu.rf_ram.memory\[71\]\[7\] _01779_ _01780_ _02508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_55_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08152__A1 _03412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08637_ _03719_ _00525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05849_ _01484_ _01486_ _01487_ _01488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06702__A2 _02313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06553__I2 u_cpu.rf_ram.memory\[138\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11387__CLK net220 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08568_ _03676_ _03668_ _03677_ _00498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout10 net11 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout21 net25 net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_23_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout32 net33 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_07519_ u_cpu.rf_ram.memory\[44\]\[6\] _02990_ _02999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout43 net50 net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_08499_ _03564_ u_cpu.rf_ram.memory\[13\]\[1\] _03633_ _03635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08455__A2 _03202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout54 net55 net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_70_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout65 net71 net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout76 net78 net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_10_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10530_ _05057_ _05061_ _05070_ _01068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06466__A1 _02078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout87 net89 net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_11_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout98 net99 net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__06561__S1 _02174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10461_ _04492_ _05019_ _04700_ _04581_ _05020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_10_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08207__A2 _03438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12200_ _00883_ net399 u_cpu.rf_ram.memory\[113\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11211__A1 _05462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10392_ _04975_ _01025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12131_ _00814_ net436 u_cpu.rf_ram.memory\[122\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12062_ _00745_ net285 u_cpu.rf_ram.memory\[35\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07718__A1 _01820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11013_ u_cpu.rf_ram.memory\[86\]\[2\] _05372_ _05373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06077__S0 _01692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09951__I _04443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[30\]_CLK net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12162__CLK net497 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06796__B _01709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07471__I _02939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11915_ _00611_ net463 u_cpu.rf_ram.memory\[130\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08694__A2 _03753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09891__A1 u_cpu.rf_ram.memory\[114\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06544__I2 u_cpu.rf_ram.memory\[70\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06087__I _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[45\]_CLK net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11846_ _00542_ net421 u_cpu.rf_ram.memory\[39\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09643__A1 u_arbiter.i_wb_cpu_rdt\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11777_ _00473_ net150 u_cpu.rf_ram.memory\[13\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10253__A2 _03123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10728_ _05187_ _05192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_13_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout123_I net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10659_ _05148_ _05133_ _05149_ _01118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09946__A2 _04572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06304__S1 _01774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12329_ _01009_ net504 u_cpu.cpu.ctrl.o_ibus_adr\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout492_I net493 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12505__CLK net168 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07870_ _03191_ _03229_ _03235_ _00242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08382__A1 _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06821_ u_cpu.rf_ram.memory\[140\]\[6\] u_cpu.rf_ram.memory\[141\]\[6\] u_cpu.rf_ram.memory\[142\]\[6\]
+ u_cpu.rf_ram.memory\[143\]\[6\] _02169_ _01816_ _02432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_42_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08509__I0 _03574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09540_ _04303_ _00845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_95_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11269__A1 _02915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06752_ _02078_ _02362_ _02363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08477__I _03620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07381__I _02903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08134__A1 u_cpu.rf_ram.memory\[62\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09471_ u_cpu.rf_ram.memory\[115\]\[6\] _04245_ _04254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06683_ u_cpu.rf_ram.memory\[44\]\[5\] u_cpu.rf_ram.memory\[45\]\[5\] u_cpu.rf_ram.memory\[46\]\[5\]
+ u_cpu.rf_ram.memory\[47\]\[5\] _01721_ _01879_ _02295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_64_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10021__B _02680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08685__A2 _03747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09882__A1 _04244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08422_ _03585_ _00444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06791__S1 _01676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08353_ u_cpu.rf_ram.memory\[53\]\[3\] _03541_ _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09634__A1 u_arbiter.i_wb_cpu_rdt\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07304_ _02845_ _02846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06448__A1 _02060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08284_ _03497_ _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07235_ u_cpu.rf_ram.memory\[21\]\[7\] _02791_ _02802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09937__A2 _04456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08940__I _02766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07166_ u_cpu.rf_ram.memory\[82\]\[1\] _02741_ _02747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06117_ _01719_ _01724_ _01727_ _01732_ _01733_ _01734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_133_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07097_ _02549_ _02681_ _02682_ _02687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_69_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06460__I _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06048_ _01397_ _01665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout200 net201 net200 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_138_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12185__CLK net390 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout211 net213 net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_47_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout222 net223 net222 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout233 net235 net233 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_43_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout244 net245 net244 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout255 net262 net255 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout266 net267 net266 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_115_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09807_ u_arbiter.i_wb_cpu_rdt\[12\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[12\]
+ _04417_ _04527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06223__I1 u_cpu.rf_ram.memory\[9\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout277 net280 net277 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_86_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout288 net289 net288 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_07999_ _03259_ _03312_ _03317_ _00289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10180__A1 _04833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout299 net304 net299 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XFILLER_46_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09738_ _02616_ _04396_ _04462_ _00884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05804__I _01450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08125__A1 u_cpu.rf_ram.memory\[62\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09669_ _04255_ _04385_ _04394_ _00883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09873__A1 _02722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11700_ _00404_ net425 u_cpu.rf_ram.memory\[55\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12680_ _01358_ net96 u_cpu.rf_ram.memory\[23\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06782__S1 _01660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11631_ _00335_ net175 u_cpu.rf_ram.memory\[62\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09625__A1 u_arbiter.i_wb_cpu_rdt\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08428__A2 _03202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11562_ _00266_ net259 u_cpu.rf_ram.memory\[75\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10513_ _05059_ _05061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_11_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06534__S1 _02033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10157__I _02776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11493_ _00197_ net105 u_cpu.rf_ram.memory\[16\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10444_ _03118_ _05004_ _05005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07939__A1 _03262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11402__CLK net217 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12528__CLK net276 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10375_ u_cpu.rf_ram.memory\[109\]\[2\] _04965_ _04966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08600__A2 _03688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12114_ _00797_ net118 u_cpu.rf_ram.memory\[11\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_scanchain_local.scan_flop\[14\] u_arbiter.i_wb_cpu_rdt\[11\] net542 u_arbiter.i_wb_cpu_dbus_dat\[8\]
+ net11 u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
X_12045_ _00728_ net495 u_cpu.cpu.mem_if.signbit vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07167__A2 _02746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11552__CLK net253 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12678__CLK net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06914__A2 _02523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09864__A1 _04518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10474__A2 _05004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06142__A3 _01758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06773__S1 _02109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout240_I net247 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11829_ _00525_ net141 u_cpu.rf_ram.memory\[14\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout338_I net395 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout505_I net506 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09856__I _04397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07020_ _02569_ _02537_ _02538_ _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_31_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07376__I _02899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08971_ _03919_ _03923_ _03932_ _00646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10016__B _04710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07922_ u_cpu.rf_ram.memory\[76\]\[6\] _03260_ _03269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09591__I _04294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07853_ _03195_ _03217_ _03224_ _00236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06905__A2 _02505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06804_ _02147_ _02414_ _02415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06461__S0 _02074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07784_ u_cpu.rf_ram.memory\[40\]\[7\] _03167_ _03178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09523_ _04285_ _04287_ _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06735_ u_cpu.rf_ram.memory\[128\]\[5\] u_cpu.rf_ram.memory\[129\]\[5\] u_cpu.rf_ram.memory\[130\]\[5\]
+ u_cpu.rf_ram.memory\[131\]\[5\] _01614_ _01616_ _02347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09855__A1 _04560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09454_ _03899_ _04242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10465__A2 _04434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06666_ _02081_ _02277_ _01970_ _02278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08405_ _03575_ _00437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06764__S1 _01633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09385_ _04199_ _00794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09607__A1 u_arbiter.i_wb_cpu_rdt\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06597_ u_cpu.rf_ram.memory\[36\]\[4\] u_cpu.rf_ram.memory\[37\]\[4\] u_cpu.rf_ram.memory\[38\]\[4\]
+ u_cpu.rf_ram.memory\[39\]\[4\] _01698_ _02109_ _02210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_36_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08336_ _03501_ _03525_ _03532_ _00411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06455__I _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11425__CLK net291 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08267_ _02738_ _03484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08830__A2 _03835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09766__I _04439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07218_ _02791_ _02792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06692__I1 u_cpu.rf_ram.memory\[109\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08198_ _03412_ _03439_ _03444_ _00361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07149_ _02730_ _02731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08594__A1 _03678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06404__B _01744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11575__CLK net340 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06190__I _01606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09791__B1 _04508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10160_ _04833_ _04811_ _04834_ _00934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_79_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10091_ _04747_ _04777_ _04778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06452__S0 _01574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09846__A1 _04425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10993_ _02762_ _05359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10456__A2 _04500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12200__CLK net399 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06755__S1 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12663_ _01342_ net87 u_cpu.rf_ram.memory\[100\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06380__I0 u_cpu.rf_ram.memory\[32\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11271__I _05534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05883__A2 _01481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11614_ _00318_ net239 u_cpu.rf_ram.memory\[64\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12594_ _01273_ net279 u_cpu.rf_ram.memory\[88\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07085__A1 _02675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11545_ _00249_ net258 u_cpu.rf_ram.memory\[74\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08821__A2 _03835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11918__CLK net457 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11476_ _00180_ net111 u_cpu.rf_ram.memory\[4\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10427_ _04808_ _04993_ _04995_ _01040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07196__I _02771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08585__A1 _03666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10358_ _02571_ _01412_ _01379_ _04952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_48_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10289_ _04912_ _00985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_97_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07924__I _03086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12028_ _00711_ net320 u_cpu.rf_ram.memory\[91\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout190_I net191 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10144__A1 _04821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout288_I net289 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06443__S0 _01826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06899__A1 _01778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10695__A2 _05168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout455_I net460 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09837__A1 _04436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06520_ u_cpu.rf_ram.memory\[112\]\[3\] u_cpu.rf_ram.memory\[113\]\[3\] u_cpu.rf_ram.memory\[114\]\[3\]
+ u_cpu.rf_ram.memory\[115\]\[3\] _02133_ _01908_ _02134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_59_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08755__I _03789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06746__S1 _02071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06451_ _01564_ _02000_ _02065_ _00002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11448__CLK net299 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09170_ _04057_ _04059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06382_ _01993_ _01995_ _01996_ _01997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_33_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08121_ _03393_ _03394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07076__A1 _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08812__A2 _03822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11598__CLK net251 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08052_ _03083_ _03351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06674__I1 u_cpu.rf_ram.memory\[49\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07003_ _02564_ _02609_ _02610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_11_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08576__A1 u_cpu.rf_ram.memory\[71\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07379__A2 _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08954_ _03921_ _03923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07905_ _03067_ _03257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10135__A1 _04814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08885_ _03875_ _00617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10686__A2 _05165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07836_ u_cpu.rf_ram.memory\[129\]\[7\] _03203_ _03214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12223__CLK net343 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07551__A2 _03020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07767_ _03167_ _03168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09506_ u_cpu.rf_ram.memory\[33\]\[3\] _04274_ _04276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06718_ _02150_ _02329_ _02153_ _02330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07698_ _03112_ _03119_ _00186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06737__S1 _02174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09437_ _04147_ _04226_ _04231_ _00814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06649_ u_cpu.rf_ram.memory\[132\]\[4\] u_cpu.rf_ram.memory\[133\]\[4\] u_cpu.rf_ram.memory\[134\]\[4\]
+ u_cpu.rf_ram.memory\[135\]\[4\] _02061_ _02174_ _02262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_125_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12373__CLK net344 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06185__I _01777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09368_ _02854_ _04188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09056__A2 _03978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07067__A1 _01430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08319_ u_cpu.rf_ram.memory\[55\]\[6\] _03517_ _03522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09299_ u_cpu.rf_ram.memory\[120\]\[0\] _04143_ _04144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08803__A2 _03822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11330_ _00034_ net68 u_cpu.rf_ram.memory\[21\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07082__A4 _02563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11261_ _02903_ _05523_ _05529_ _01340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08567__A1 u_cpu.rf_ram.memory\[71\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10212_ _04864_ _00956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11192_ _05098_ _03165_ _05488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10143_ u_cpu.rf_ram.memory\[32\]\[3\] _04818_ _04822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06788__C _01606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10074_ _04602_ _04642_ _04553_ _04609_ _04762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_94_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[7\] u_arbiter.i_wb_cpu_rdt\[4\] net548 u_arbiter.i_wb_cpu_dbus_dat\[1\]
+ net15 u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_47_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10677__A2 _05152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07542__A2 _03011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09819__A1 _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08575__I _03506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10429__A2 _04993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10976_ _05286_ _05337_ _05346_ _01238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05856__A2 _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12646_ _01325_ net123 u_cpu.rf_ram.memory\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09047__A2 _03978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06105__I0 u_cpu.rf_ram.memory\[104\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12577_ _01256_ net168 u_cpu.rf_ram.memory\[111\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11528_ _00232_ net511 u_cpu.rf_ram.memory\[139\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06900__S1 _01763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10345__I _04908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout203_I net208 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06281__A2 _01896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11459_ _00163_ net222 u_cpu.rf_ram.memory\[47\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08558__A1 _03666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10365__A1 _02700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07230__A1 _02763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05951_ _01567_ _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10117__A1 _04532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08670_ u_cpu.rf_ram.memory\[39\]\[3\] _03738_ _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05882_ u_cpu.cpu.ctrl.o_ibus_adr\[17\] _01511_ _01514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_27_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10013__C _04503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06187__I3 u_cpu.rf_ram.memory\[79\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07533__A2 _03008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07621_ _03060_ _03064_ _03066_ _00162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_19_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07552_ _03021_ _03022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09286__A2 _04129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06503_ _01665_ _02117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07297__A1 _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07483_ _02900_ _02969_ _02974_ _00116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06434_ _01802_ _02048_ _01805_ _02049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09222_ _04092_ _04097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10840__A2 _05261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09153_ _03975_ _04045_ _04048_ _00712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06365_ _01656_ _01979_ _01867_ _01980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_120_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08104_ _03335_ _03382_ _03384_ _00327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08797__A1 _03819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06647__I1 u_cpu.rf_ram.memory\[129\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09084_ u_cpu.rf_ram.memory\[37\]\[0\] _04004_ _04005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06296_ _01751_ _01911_ _01755_ _01912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_120_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08035_ _03335_ _03337_ _03339_ _00303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06272__A2 _01875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08549__A1 u_cpu.rf_ram.memory\[73\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10356__A1 u_cpu.cpu.ctrl.o_ibus_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10191__S _04849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07221__A1 _02740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09986_ _04494_ _04679_ _04681_ _04683_ _04684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_66_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07772__A2 _03168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08937_ _03909_ _03910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11613__CLK net238 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06407__S0 _01752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10659__A2 _05133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08868_ _03824_ _03859_ _03865_ _00610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08721__A1 _03757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07819_ _03203_ _03204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08799_ _03815_ _03822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10830_ _04091_ _03310_ _05256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11763__CLK net491 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07288__A1 _02746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10761_ u_cpu.rf_ram.memory\[79\]\[5\] _05207_ _05214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10292__B1 _04910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12500_ _01179_ net37 u_cpu.rf_ram.memory\[107\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05838__A2 _01461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10692_ _05140_ _05164_ _05170_ _01130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09029__A2 _03959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12431_ _01110_ net358 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09985__B1 _04682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12362_ _01041_ net211 u_cpu.rf_ram.memory\[93\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10595__A1 u_cpu.rf_ram.memory\[28\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11313_ _02648_ _02650_ u_cpu.rf_ram.rdata\[7\] _05560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__07460__A1 _02900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12293_ _00975_ net496 u_cpu.cpu.bufreg.lsb\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_101_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[5\]_D u_arbiter.i_wb_cpu_rdt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12269__CLK net530 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07675__S _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11244_ u_cpu.rf_ram.memory\[98\]\[5\] _05515_ _05519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11175_ u_cpu.rf_ram.memory\[25\]\[0\] _05478_ _05479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10126_ _04807_ _04808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07763__A2 _03155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05774__A1 u_cpu.cpu.immdec.imm24_20\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10057_ _04542_ _04745_ _04746_ _00919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_23_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08712__A1 _03745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07279__A1 _01658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout153_I net154 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10959_ _05335_ _05337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10822__A2 _05249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout320_I net322 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12629_ _01308_ net53 u_cpu.rf_ram.memory\[25\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08779__A1 _03755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06150_ _01704_ _01767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_106_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10586__A1 _05046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09440__A2 _04230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06081_ _01650_ _01698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__07451__A1 _02921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10008__C _04555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09840_ _04499_ _04543_ _04556_ _04557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10889__A2 _05289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07384__I _02762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06502__B _02115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08951__A1 _03919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07754__A2 _03158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09771_ _03118_ _04493_ _04494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06983_ _01412_ _02589_ _02590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08722_ u_cpu.rf_ram.memory\[49\]\[5\] _03770_ _03774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05934_ u_cpu.cpu.ctrl.o_ibus_adr\[28\] _01547_ _01548_ _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_6_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout66_I net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11786__CLK net350 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08703__A1 u_cpu.rf_ram.memory\[137\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05865_ _01489_ _01498_ _01499_ _01500_ u_arbiter.o_wb_cpu_adr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_08653_ _03678_ _03722_ _03729_ _00531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10510__A1 _05057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07604_ _02992_ _03048_ _03054_ _00157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05796_ _01442_ _01443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_81_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08584_ u_cpu.rf_ram.memory\[70\]\[0\] _03688_ _03689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07535_ _03006_ _03011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10813__A2 _05246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06868__I1 u_cpu.rf_ram.memory\[109\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07466_ _02910_ _02955_ _02962_ _00111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09205_ _02585_ _02586_ _02553_ _02559_ _04085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_91_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06417_ _01766_ _02030_ _02031_ _02032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_33_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07397_ _02915_ _02916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09136_ net2 _04026_ _04037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06348_ _01597_ _01962_ _01603_ _01963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12411__CLK net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09431__A2 _04227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10577__A1 _05098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09067_ _03975_ _03991_ _03994_ _00680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07442__A1 _02904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06279_ _01667_ _01895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_120_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09774__I _04426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08018_ u_cpu.rf_ram.memory\[66\]\[2\] _03328_ _03329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07993__A2 _03313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09195__A1 _02673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12561__CLK net162 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09969_ _01443_ u_arbiter.i_wb_cpu_rdt\[9\] _04669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[11\]_SE net544 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11931_ _00627_ net419 u_cpu.rf_ram.memory\[22\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10501__A1 _05051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11862_ _00558_ net420 u_cpu.rf_ram.memory\[49\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09014__I _03957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10813_ u_cpu.rf_ram.memory\[107\]\[0\] _05246_ _05247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11793_ _00489_ net352 u_cpu.rf_ram.memory\[73\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11509__CLK net301 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10744_ _05200_ _05202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10804__A2 _05233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10675_ _05144_ _05152_ _05159_ _01124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12091__CLK net403 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12414_ _01093_ net82 u_cpu.rf_ram.memory\[28\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06373__I _01609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10568__A1 _05055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10109__B _04526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11659__CLK net182 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[44\] u_scanchain_local.module_data_in\[43\] net559 u_arbiter.o_wb_cpu_adr\[6\]
+ net27 u_scanchain_local.module_data_in\[44\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
X_12345_ _01024_ net112 u_cpu.rf_ram.memory\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07984__A2 _03300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12276_ _00959_ net533 u_arbiter.i_wb_cpu_dbus_adr\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11227_ _05508_ _01327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06619__S0 _02136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07736__A2 _03146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11158_ _05449_ _05465_ _05468_ _01298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10740__A1 _05148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10109_ _01442_ u_arbiter.i_wb_cpu_rdt\[19\] _04526_ _04793_ _04794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_11089_ _02693_ _01393_ _05419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09489__A2 _04258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout270_I net271 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11296__A2 _05547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout368_I net372 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08161__A2 _03408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[38\]_D u_scanchain_local.module_data_in\[37\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11048__A2 _05393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout535_I net536 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output7_I net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07320_ _02859_ _00068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09110__A1 _03977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09661__A2 _04384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07251_ u_cpu.rf_ram.memory\[81\]\[4\] _02810_ _02813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06202_ _01568_ _01819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07182_ _02748_ u_cpu.rf_ram_if.wdata1_r\[4\] _02760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_9_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10559__A1 u_cpu.rf_ram.memory\[96\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06133_ _01746_ _01749_ _01750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06227__A2 _01842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12584__CLK net207 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07975__A2 _03299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06064_ _01426_ _01681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10533__I _05071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout404 net407 net404 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout415 net417 net415 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA_u_scanchain_local.scan_flop\[34\]_SE net549 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout426 net429 net426 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__07727__A2 _03143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09823_ _04485_ _04438_ _04525_ _04540_ _04541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
Xfanout437 net442 net437 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout448 net449 net448 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06786__I0 u_cpu.rf_ram.memory\[96\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout459 net460 net459 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10731__A1 u_cpu.rf_ram.memory\[99\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09754_ _04475_ _04477_ _04478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06250__I2 u_cpu.rf_ram.memory\[50\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06966_ _02568_ _02565_ _02570_ _02573_ _02574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_80_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08705_ _03509_ _03763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05917_ _01537_ _01535_ _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09685_ _01440_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[12\] _04410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__06538__I0 u_cpu.rf_ram.memory\[84\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06897_ _01797_ _02506_ _02507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08152__A2 _03407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08636_ _03574_ u_cpu.rf_ram.memory\[14\]\[6\] _03711_ _03719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[29\]_D u_arbiter.i_wb_cpu_rdt\[26\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_05848_ _01484_ _01486_ _01455_ _01487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11039__A2 _05384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08567_ u_cpu.rf_ram.memory\[71\]\[3\] _03674_ _03677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05779_ _01400_ _01429_ _00025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xfanout11 net14 net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09101__A1 _02830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout22 net24 net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout33 net34 net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_07518_ _02912_ _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout44 net45 net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_126_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08498_ _03634_ _00471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10798__A1 _05206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout55 net62 net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout66 net71 net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout77 net78 net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__06466__A2 _02079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07663__A1 u_cpu.rf_ram.memory\[50\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10708__I _05175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout88 net89 net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_07449_ u_cpu.rf_ram.memory\[42\]\[7\] _02941_ _02952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11801__CLK net368 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout99 net100 net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_7_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07289__I _02832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10460_ _04401_ _04520_ _05019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06193__I _01404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09119_ u_cpu.rf_ram.memory\[36\]\[7\] _04014_ _04025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07415__A1 _02900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10391_ _04188_ u_cpu.rf_ram.memory\[3\]\[1\] _04973_ _04975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12130_ _00813_ net405 u_cpu.rf_ram.memory\[122\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06921__I _02529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05977__A1 _01590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10970__A1 _05280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09168__A1 _02731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08215__I0 _02858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12061_ _00744_ net307 u_cpu.rf_ram.memory\[35\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07953__S _03289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08915__A1 _03832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11012_ _05367_ _05372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06077__S1 _01693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12307__CLK net492 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06529__I0 u_cpu.rf_ram.memory\[92\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09340__A1 _04156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11914_ _00610_ net469 u_cpu.rf_ram.memory\[130\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06154__A1 _01766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11331__CLK net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12457__CLK net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10111__C _04795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06544__I3 u_cpu.rf_ram.memory\[71\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11845_ _00541_ net432 u_cpu.rf_ram.memory\[39\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09679__I _03114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11776_ _00472_ net149 u_cpu.rf_ram.memory\[13\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10789__A1 _02937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10727_ _05135_ _05188_ _05191_ _01144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11481__CLK net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07654__A1 u_cpu.rf_ram.memory\[50\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10658_ u_cpu.rf_ram.memory\[101\]\[7\] _05131_ _05149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07406__A1 _02921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11202__A2 _05493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout116_I net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10589_ u_cpu.rf_ram.memory\[28\]\[4\] _05104_ _05107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07927__I _02922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[57\]_SE net562 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12328_ _01008_ net504 u_cpu.cpu.ctrl.o_ibus_adr\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09159__A1 u_cpu.rf_ram.memory\[91\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10961__A1 _05268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12259_ _00942_ net90 u_cpu.rf_ram.memory\[31\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08906__A1 u_cpu.rf_ram.memory\[22\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout485_I net487 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08382__A2 _03550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06820_ _01825_ _02430_ _02431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11269__A2 _05524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06751_ u_cpu.rf_ram.memory\[20\]\[6\] u_cpu.rf_ram.memory\[21\]\[6\] u_cpu.rf_ram.memory\[22\]\[6\]
+ u_cpu.rf_ram.memory\[23\]\[6\] _01631_ _01965_ _02362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_77_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09331__A1 u_cpu.rf_ram.memory\[118\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09470_ _03915_ _04253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06682_ _01876_ _02293_ _02294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08421_ _03572_ u_cpu.rf_ram.memory\[15\]\[5\] _03578_ _03585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_52_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09619__C1 _04327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11824__CLK net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08352_ _03494_ _03537_ _03542_ _00417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout29_I net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07303_ u_cpu.rf_ram_if.wdata0_r\[0\] u_cpu.rf_ram_if.wdata1_r\[0\] _02844_ _02845_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07645__A1 u_cpu.rf_ram.memory\[47\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06448__A2 _02062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08283_ _02756_ _03497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06227__B _01588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07234_ _02773_ _02793_ _02801_ _00040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07165_ _02745_ _02746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06116_ _01605_ _01733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08070__A1 u_cpu.rf_ram.memory\[64\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07096_ _02684_ _02586_ _02685_ _02686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_69_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06047_ _01656_ _01661_ _01663_ _01664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout201 net202 net201 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_120_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout212 net213 net212 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout223 net229 net223 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout234 net235 net234 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__10704__A1 u_cpu.rf_ram.memory\[104\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout245 net246 net245 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_43_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout256 net257 net256 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_09806_ _04446_ _04526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout267 net268 net267 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_75_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08373__A2 _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout278 net279 net278 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__11354__CLK net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07998_ u_cpu.rf_ram.memory\[67\]\[2\] _03316_ _03317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07572__I _03033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10180__A2 _04837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout289 net290 net289 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09737_ _04398_ _04461_ _04462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06949_ _01372_ _02557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_55_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09322__A1 _04158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08125__A2 _03395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06188__I _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09668_ u_cpu.rf_ram.memory\[113\]\[7\] _04383_ _04394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09873__A2 _04224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08619_ _03682_ _03701_ _03709_ _00517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07884__A1 u_cpu.rf_ram.memory\[74\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09599_ _04349_ _00858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11630_ _00334_ net181 u_cpu.rf_ram.memory\[63\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09625__A2 _04293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11561_ _00265_ net258 u_cpu.rf_ram.memory\[75\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10512_ _05059_ _05060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11492_ _00196_ net105 u_cpu.rf_ram.memory\[16\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10443_ _02674_ _02704_ _05004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11196__A1 _05444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10243__I0 u_arbiter.i_wb_cpu_dbus_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07939__A2 _03274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08061__A1 u_cpu.rf_ram.memory\[64\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10374_ _04960_ _04965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12113_ _00796_ net125 u_cpu.rf_ram.memory\[11\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06611__A2 _02223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07683__S _03101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09936__I0 u_arbiter.i_wb_cpu_rdt\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12044_ _00727_ net480 u_cpu.cpu.state.genblk1.misalign_trap_sync_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_78_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08578__I _03509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10171__A2 _04840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11847__CLK net508 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09313__A1 _04152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08116__A2 _03386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10459__B1 _04491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06098__I _01665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11120__A1 u_cpu.cpu.ctrl.i_iscomp vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09403__S _04202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06517__I3 u_cpu.rf_ram.memory\[123\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11828_ _00524_ net144 u_cpu.rf_ram.memory\[14\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11997__CLK net400 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09616__A2 _04352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout233_I net235 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11759_ _00455_ net479 u_cpu.rf_ram.memory\[141\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06047__B _01663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout400_I net402 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11187__A1 _05458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10934__A1 _05282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11179__I _05476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08970_ u_cpu.rf_ram.memory\[127\]\[7\] _03921_ _03932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11377__CLK net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07921_ _03083_ _03268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12622__CLK net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08355__A2 _03541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10811__I _05244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07852_ u_cpu.rf_ram.memory\[139\]\[5\] _03220_ _03224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07392__I _02772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06803_ u_cpu.rf_ram.memory\[80\]\[6\] u_cpu.rf_ram.memory\[81\]\[6\] u_cpu.rf_ram.memory\[82\]\[6\]
+ u_cpu.rf_ram.memory\[83\]\[6\] _01651_ _02033_ _02414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_84_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput1 io_in[0] net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_56_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06461__S1 _01599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07783_ _03084_ _03169_ _03177_ _00213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09522_ _03125_ _04286_ _04287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06734_ _01830_ _02345_ _01628_ _02346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06937__S u_arbiter.i_wb_cpu_dbus_we vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11111__A1 u_cpu.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09855__A2 _04562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09453_ _04237_ _04239_ _04241_ _00820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06665_ u_cpu.rf_ram.memory\[16\]\[5\] u_cpu.rf_ram.memory\[17\]\[5\] u_cpu.rf_ram.memory\[18\]\[5\]
+ u_cpu.rf_ram.memory\[19\]\[5\] _01852_ _01968_ _02277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_25_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08404_ _03574_ u_cpu.rf_ram.memory\[9\]\[6\] _03561_ _03575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09384_ _04198_ u_cpu.rf_ram.memory\[8\]\[6\] _04185_ _04199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_24_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12002__CLK net415 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09607__A2 _04326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06596_ _01988_ _02208_ _02107_ _02209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_33_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08335_ u_cpu.rf_ram.memory\[54\]\[4\] _03529_ _03532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08266_ _03423_ _03474_ _03483_ _00390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12152__CLK net398 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07217_ _02786_ _02790_ _02791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11178__A1 _05449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08197_ u_cpu.rf_ram.memory\[19\]\[2\] _03443_ _03444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07148_ _02701_ _02725_ _02729_ _02730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_133_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10925__A1 _05273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09791__A1 _02633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07079_ _02556_ _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09782__I _04399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[44\]_CLK net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10090_ _04550_ _04700_ _04777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09543__A1 _04285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08346__A2 _03538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06452__S1 _01838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[59\]_CLK net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11102__A1 _01382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10992_ _05357_ _05349_ _05358_ _01242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09846__A2 _04561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07857__A1 _03199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12662_ _01341_ net159 u_cpu.rf_ram.memory\[100\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06380__I1 u_cpu.rf_ram.memory\[33\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11613_ _00317_ net238 u_cpu.rf_ram.memory\[64\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12593_ _01272_ net278 u_cpu.rf_ram.memory\[88\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07085__A2 _02676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11544_ _00248_ net261 u_cpu.rf_ram.memory\[74\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08282__A1 _03494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11475_ _00179_ net121 u_cpu.rf_ram.memory\[4\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06683__I2 u_cpu.rf_ram.memory\[46\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11169__A1 _05460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09893__S _01441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06381__I _01662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10426_ u_cpu.rf_ram.memory\[93\]\[0\] _04994_ _04995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12645__CLK net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10916__A1 _05284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10357_ _04951_ _01014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_125_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10288_ u_arbiter.i_wb_cpu_ibus_adr\[1\] _04907_ _04910_ _01444_ _04912_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_111_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08337__A2 _03529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12027_ _00710_ net492 u_cpu.cpu.state.o_cnt_r\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06348__A1 _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06330__B _01823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05725__I u_cpu.cpu.branch_op vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06443__S1 _01827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout183_I net184 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12025__CLK net490 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09837__A2 _04523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout350_I net354 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout448_I net449 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06450_ _02053_ _02064_ _02065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06371__I1 u_cpu.rf_ram.memory\[41\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12175__CLK net386 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06381_ _01662_ _01996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10455__I0 u_cpu.cpu.immdec.imm11_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08120_ _02920_ _03005_ _03393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07076__A2 _02658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08273__A1 _03485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08051_ _03349_ _03338_ _03350_ _00308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_70_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06674__I2 u_cpu.rf_ram.memory\[50\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07002_ _02607_ u_cpu.cpu.ctrl.i_iscomp _02608_ _02609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08025__A1 _03266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10907__A1 u_cpu.rf_ram.memory\[84\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09773__A1 _04484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08576__A2 _03674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09816__B _04532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10383__A2 _04965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout96_I net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08953_ _03921_ _03922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08328__A2 _03526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07904_ _03252_ _03254_ _03256_ _00255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08884_ _03566_ u_cpu.rf_ram.memory\[12\]\[2\] _03872_ _03875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07835_ _03197_ _03205_ _03213_ _00229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07766_ _03018_ _03166_ _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09505_ _04244_ _04270_ _04275_ _00838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06717_ u_cpu.rf_ram.memory\[84\]\[5\] u_cpu.rf_ram.memory\[85\]\[5\] u_cpu.rf_ram.memory\[86\]\[5\]
+ u_cpu.rf_ram.memory\[87\]\[5\] _01922_ _02151_ _02329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10189__S _04849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07697_ u_cpu.cpu.state.genblk1.misalign_trap_sync_r u_cpu.cpu.state.stage_two_req
+ _03118_ _03119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_72_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12518__CLK net203 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09436_ u_cpu.rf_ram.memory\[122\]\[2\] _04230_ _04231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08882__S _03872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06648_ _01947_ _02260_ _02261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_55_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09367_ _04187_ _00788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06579_ u_cpu.rf_ram.memory\[28\]\[4\] u_cpu.rf_ram.memory\[29\]\[4\] u_cpu.rf_ram.memory\[30\]\[4\]
+ u_cpu.rf_ram.memory\[31\]\[4\] _02084_ _01577_ _02192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_90_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08318_ _03504_ _03514_ _03521_ _00404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11542__CLK net250 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08264__A1 _03421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12668__CLK net286 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09298_ _04141_ _04143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_123_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10071__A1 _01391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08249_ _03472_ _03474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06665__I2 u_cpu.rf_ram.memory\[18\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08016__A1 _03257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11260_ u_cpu.rf_ram.memory\[100\]\[3\] _05527_ _05529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09764__A1 _04429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10211_ u_arbiter.i_wb_cpu_dbus_adr\[15\] u_arbiter.i_wb_cpu_dbus_adr\[14\] _04861_
+ _04864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08567__A2 _03674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11191_ _05462_ _05478_ _05487_ _01312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10142_ _04820_ _04821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09516__A1 u_cpu.cpu.bufreg.lsb\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08319__A2 _03517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10073_ _04652_ _04760_ _04761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12048__CLK net379 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07961__S _03289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09819__A2 _04396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10975_ u_cpu.rf_ram.memory\[85\]\[7\] _05335_ _05346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_95_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12645_ _01324_ net124 u_cpu.rf_ram.memory\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12576_ _01255_ net168 u_cpu.rf_ram.memory\[111\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11527_ _00231_ net488 u_cpu.rf_ram.memory\[139\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06325__B _01810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08007__A1 _03268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11458_ _00162_ net222 u_cpu.rf_ram.memory\[47\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07000__I u_cpu.cpu.state.o_cnt_r\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09755__A1 _04474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10409_ _04188_ u_cpu.rf_ram.memory\[2\]\[1\] _04983_ _04985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06113__S0 _01729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11389_ _00093_ net182 u_cpu.rf_ram.memory\[78\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07230__A2 _02792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout398_I net399 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09507__A1 _04247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05950_ _01390_ _01392_ _01396_ _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_87_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10117__A2 _04710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05881_ _01505_ _01510_ _01511_ _01513_ u_arbiter.o_wb_cpu_adr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA_fanout565_I net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11415__CLK net224 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07620_ u_cpu.rf_ram.memory\[47\]\[0\] _03065_ _03066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06741__A1 _01406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07551_ _03018_ _03020_ _03021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06502_ _01566_ _02077_ _02089_ _02115_ _02116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11565__CLK net341 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08494__A1 _03606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07482_ u_cpu.rf_ram.memory\[45\]\[2\] _02973_ _02974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09221_ _04061_ _04093_ _04096_ _00733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06433_ u_cpu.rf_ram.memory\[76\]\[2\] u_cpu.rf_ram.memory\[77\]\[2\] u_cpu.rf_ram.memory\[78\]\[2\]
+ u_cpu.rf_ram.memory\[79\]\[2\] _02047_ _01803_ _02048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_61_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout11_I net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09152_ u_cpu.rf_ram.memory\[91\]\[1\] _04046_ _04048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08246__A1 _03423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06364_ u_cpu.rf_ram.memory\[48\]\[2\] u_cpu.rf_ram.memory\[49\]\[2\] u_cpu.rf_ram.memory\[50\]\[2\]
+ u_cpu.rf_ram.memory\[51\]\[2\] _01657_ _01660_ _01979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08103_ u_cpu.rf_ram.memory\[63\]\[0\] _03383_ _03384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09994__A1 _01440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08797__A2 _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06295_ u_cpu.rf_ram.memory\[116\]\[1\] u_cpu.rf_ram.memory\[117\]\[1\] u_cpu.rf_ram.memory\[118\]\[1\]
+ u_cpu.rf_ram.memory\[119\]\[1\] _01752_ _01753_ _01911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09083_ _04002_ _04004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_11_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08034_ u_cpu.rf_ram.memory\[65\]\[0\] _03338_ _03339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08549__A2 _03659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10356__A2 _04906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07845__I _03215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10600__I0 u_arbiter.i_wb_cpu_rdt\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07221__A2 _02792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09985_ _04680_ _04609_ _04682_ _04652_ _04575_ _04683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_118_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08936_ _02761_ _03909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10108__A2 _04310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11305__A1 _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06980__A1 _02553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08867_ u_cpu.rf_ram.memory\[130\]\[3\] _03863_ _03865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07818_ _02804_ _03202_ _03203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08798_ _03493_ _03821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11908__CLK net461 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07749_ u_cpu.rf_ram.memory\[17\]\[1\] _03155_ _03157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06196__I _01812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10760_ _04826_ _05213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07288__A2 _02833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09419_ u_cpu.rf_ram.memory\[112\]\[4\] _04217_ _04220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10691_ u_cpu.rf_ram.memory\[103\]\[3\] _05168_ _05170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12430_ _01109_ net363 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10044__A1 _02529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09985__A1 _04680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12361_ _01040_ net211 u_cpu.rf_ram.memory\[93\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09985__B2 _04652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10595__A2 _05099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11312_ _04907_ _05558_ _05559_ _01361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_10_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12292_ _00974_ net495 u_cpu.cpu.bufreg.lsb\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07460__A2 _02954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09737__A1 _04398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11243_ _05456_ _05511_ _05518_ _01333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11174_ _05476_ _05478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_49_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11277__I _05534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08960__A2 _03926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10125_ _02738_ _04807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06810__I2 u_cpu.rf_ram.memory\[70\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05774__A2 _01389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[8\]_SE net549 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10056_ u_cpu.cpu.csr_imm _02530_ _04482_ _04736_ _04746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_76_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07279__A2 _02719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10958_ _05335_ _05336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_16_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10283__A1 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout146_I net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10889_ _05278_ _05289_ _05295_ _01202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12628_ _01307_ net53 u_cpu.rf_ram.memory\[25\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10035__A1 _04416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09976__A1 u_cpu.cpu.immdec.imm30_25\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08779__A2 _03802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06629__I2 u_cpu.rf_ram.memory\[86\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout313_I net314 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12559_ _01238_ net213 u_cpu.rf_ram.memory\[85\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06334__S0 _01831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12213__CLK net318 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06080_ _01648_ _01697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07451__A2 _02940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09728__A1 _04439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10338__A2 _04936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12363__CLK net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09770_ _04438_ _04445_ _04493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08951__A2 _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06982_ _02588_ _02533_ _02546_ _02589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_101_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06962__A1 _02569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05765__A2 _01388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08721_ _03757_ _03766_ _03773_ _00555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05933_ _01489_ _01552_ _01553_ u_arbiter.o_wb_cpu_adr\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08703__A2 _03753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08496__I _03632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08652_ u_cpu.rf_ram.memory\[138\]\[4\] _03726_ _03729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05864_ u_arbiter.i_wb_cpu_dbus_adr\[13\] _01493_ _01500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06714__A1 _01740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout59_I net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10510__A2 _05042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07603_ u_cpu.rf_ram.memory\[48\]\[3\] _03052_ _03054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08583_ _03686_ _03688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05795_ _01441_ _01442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_39_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07534_ _02987_ _03007_ _03010_ _00131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07465_ u_cpu.rf_ram.memory\[46\]\[5\] _02958_ _02962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09204_ _01409_ _02556_ _04080_ _04082_ _04084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_22_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06416_ _01678_ _02031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07396_ _02777_ _02915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10026__A1 _01440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09135_ _03112_ _04036_ _00706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06347_ u_cpu.rf_ram.memory\[0\]\[2\] u_cpu.rf_ram.memory\[1\]\[2\] u_cpu.rf_ram.memory\[2\]\[2\]
+ u_cpu.rf_ram.memory\[3\]\[2\] _01598_ _01599_ _01962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_108_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10577__A2 _02982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09066_ u_cpu.rf_ram.memory\[38\]\[1\] _03992_ _03994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06278_ _01720_ _01893_ _01723_ _01894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07442__A2 _02942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09719__A1 _04437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08017_ _03323_ _03328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12706__CLK net353 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09195__A2 _02677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06253__I0 u_cpu.rf_ram.memory\[60\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08942__A2 _03904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09968_ _03115_ u_arbiter.i_wb_cpu_rdt\[25\] _04668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05756__A2 u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08919_ _03895_ _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_44_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09899_ _04549_ _04455_ _04604_ _04605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11930_ _00626_ net419 u_cpu.rf_ram.memory\[22\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06919__I _02527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11861_ _00557_ net377 u_cpu.rf_ram.memory\[49\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10812_ _05244_ _05246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11792_ _00488_ net373 u_cpu.rf_ram.memory\[73\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10743_ _05200_ _05201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_40_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12236__CLK net264 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10674_ u_cpu.rf_ram.memory\[102\]\[5\] _05155_ _05159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12413_ _01092_ net90 u_cpu.rf_ram.memory\[28\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12344_ _00021_ net385 u_cpu.cpu.alu.add_cy_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_scanchain_local.scan_flop\[37\] u_scanchain_local.module_data_in\[36\] net556 u_arbiter.i_wb_cpu_dbus_dat\[31\]
+ net24 u_scanchain_local.module_data_in\[37\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
X_12275_ _00958_ net533 u_arbiter.i_wb_cpu_dbus_adr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06603__B _02215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11226_ _02869_ u_cpu.rf_ram.memory\[0\]\[6\] _05500_ _05508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09914__B _04619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11157_ u_cpu.rf_ram.memory\[26\]\[1\] _05466_ _05468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06944__A1 _02530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06795__I1 u_cpu.rf_ram.memory\[117\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10108_ _01442_ _04310_ _04793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11088_ _05417_ _05418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10039_ _02674_ _02625_ _04466_ _04733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout263_I net264 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10256__A1 u_arbiter.i_wb_cpu_dbus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout528_I net530 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07121__A1 _01394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07250_ _02758_ _02806_ _02812_ _00045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06201_ _01400_ _01817_ _01818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_121_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11603__CLK net243 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07181_ _02733_ _02758_ _02759_ _00029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06307__S0 _01922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10559__A2 _05088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06132_ u_cpu.rf_ram.memory\[112\]\[0\] u_cpu.rf_ram.memory\[113\]\[0\] u_cpu.rf_ram.memory\[114\]\[0\]
+ u_cpu.rf_ram.memory\[115\]\[0\] _01747_ _01748_ _01749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08621__A1 _03684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06063_ _01672_ _01677_ _01679_ _01680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_47_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06513__B _01731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11753__CLK net481 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10035__B _04728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07188__A1 _02748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout405 net406 net405 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_28_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06232__C _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout416 net417 net416 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_113_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09822_ _04497_ _04457_ _04503_ _04539_ _04532_ _04540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
Xfanout427 net428 net427 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout438 net440 net438 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_58_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05738__A2 _01378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout449 net475 net449 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_115_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09753_ _04476_ _04477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_101_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06965_ _02528_ _02572_ _02573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08704_ _03761_ _03748_ _03762_ _00549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05916_ _01524_ _01538_ _01540_ u_arbiter.o_wb_cpu_adr\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09684_ _04408_ _04409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_95_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08688__A1 _03750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06896_ u_cpu.rf_ram.memory\[64\]\[7\] u_cpu.rf_ram.memory\[65\]\[7\] u_cpu.rf_ram.memory\[66\]\[7\]
+ u_cpu.rf_ram.memory\[67\]\[7\] _01798_ _01799_ _02506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08635_ _03718_ _00524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10495__A1 _05046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05847_ _01485_ _01477_ _01486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_54_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08566_ _03497_ _03676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_74_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08954__I _03921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12259__CLK net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09637__B1 _04359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05778_ _01406_ _01419_ _01423_ _01428_ _01429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__05910__A2 _01512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout12 net14 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09101__A2 _02940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07517_ _02996_ _02985_ _02997_ _00127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout23 net24 net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_126_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08497_ _03560_ u_cpu.rf_ram.memory\[13\]\[0\] _03633_ _03634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_74_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout34 net35 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__06546__S0 _01934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout45 net49 net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_70_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10798__A2 _05232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout56 net58 net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout67 net70 net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__08890__S _03871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07448_ _02913_ _02943_ _02951_ _00104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout78 net84 net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_50_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout89 net91 net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_52_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07379_ _02900_ _02893_ _02902_ _00084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09118_ _03986_ _04016_ _04024_ _00701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10390_ _04974_ _01024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07415__A2 _02925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09049_ _03909_ _03982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_2_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05977__A2 _01593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10970__A2 _05336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09168__A2 _02938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12060_ _00743_ net307 u_cpu.rf_ram.memory\[35\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11011_ _05352_ _05368_ _05371_ _01248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08915__A2 _03883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08679__A1 _03684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11913_ _00609_ net469 u_cpu.rf_ram.memory\[130\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08864__I _03858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11844_ _00540_ net421 u_cpu.rf_ram.memory\[39\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09628__B1 _04319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11775_ _00471_ net137 u_cpu.rf_ram.memory\[13\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07103__A1 _01431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10789__A2 _05162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10726_ u_cpu.rf_ram.memory\[99\]\[1\] _05189_ _05191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10657_ _04832_ _05148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11776__CLK net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07406__A2 _02923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10588_ _05049_ _05100_ _05106_ _01090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06465__I0 u_cpu.rf_ram.memory\[20\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12327_ _01007_ net525 u_cpu.cpu.ctrl.o_ibus_adr\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10634__I _05131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout109_I net158 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10961__A2 _05336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09159__A2 _04049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12258_ _00941_ net79 u_cpu.rf_ram.memory\[31\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11209_ _05460_ _05490_ _05498_ _01319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08906__A2 _03886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12189_ _00872_ net497 u_arbiter.i_wb_cpu_dbus_dat\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06917__A1 _01406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07965__I0 _02870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout380_I net381 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout478_I net484 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07590__A1 _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06750_ _02354_ _02356_ _02358_ _02360_ _01807_ _02361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_77_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12401__CLK net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10477__A1 _04545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09331__A2 _04165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06681_ u_cpu.rf_ram.memory\[40\]\[5\] u_cpu.rf_ram.memory\[41\]\[5\] u_cpu.rf_ram.memory\[42\]\[5\]
+ u_cpu.rf_ram.memory\[43\]\[5\] _01736_ _02103_ _02293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_63_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07342__A1 _02784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08420_ _03584_ _00443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09619__B1 _04321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07893__A2 _03245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08351_ u_cpu.rf_ram.memory\[53\]\[2\] _03541_ _03542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10809__I _04958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07302_ _02736_ _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08282_ _03494_ _03487_ _03496_ _00393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07645__A2 _03072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07233_ u_cpu.rf_ram.memory\[21\]\[6\] _02796_ _02801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09819__B _04537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07164_ _02744_ _02745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08215__S _03451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06115_ _01728_ _01730_ _01731_ _01732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07095_ _02680_ _02614_ _02685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06046_ _01662_ _01663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_47_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout202 net209 net202 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_132_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout213 net214 net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_134_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08949__I _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout224 net228 net224 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout235 net240 net235 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_43_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout246 net247 net246 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__10704__A2 _05177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09805_ _04473_ _04525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout257 net260 net257 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout268 net269 net268 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_07997_ _03311_ _03316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout279 net280 net279 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_47_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06948_ _01371_ _02556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_09736_ _04412_ _04435_ _04448_ _04460_ _04461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_21_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12081__CLK net410 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10468__A1 _02700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09322__A2 _04143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10468__B2 _04516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09667_ _04253_ _04385_ _04393_ _00882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06879_ u_cpu.rf_ram.memory\[120\]\[7\] u_cpu.rf_ram.memory\[121\]\[7\] u_cpu.rf_ram.memory\[122\]\[7\]
+ u_cpu.rf_ram.memory\[123\]\[7\] _01674_ _01676_ _02489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_28_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08618_ u_cpu.rf_ram.memory\[143\]\[6\] _03704_ _03709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09598_ u_arbiter.i_wb_cpu_rdt\[14\] _04326_ _04321_ u_arbiter.i_wb_cpu_dbus_dat\[14\]
+ _04327_ u_arbiter.i_wb_cpu_dbus_dat\[15\] _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__07884__A2 _03242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05895__A1 _01473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08549_ u_cpu.rf_ram.memory\[73\]\[6\] _03659_ _03664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09086__A1 u_cpu.rf_ram.memory\[37\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11560_ _00264_ net258 u_cpu.rf_ram.memory\[75\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11799__CLK net368 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10511_ _04091_ _02921_ _05059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10640__A1 _05135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11491_ _00195_ net180 u_cpu.rf_ram.memory\[16\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09389__A2 _03034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10442_ _04833_ _04994_ _05003_ _01047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10373_ _04814_ _04961_ _04964_ _01017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12112_ _00795_ net137 u_cpu.rf_ram.memory\[8\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12043_ _00726_ net308 u_cpu.rf_ram.memory\[90\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09936__I1 u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08859__I _03858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12424__CLK net357 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06375__A2 _01989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06379__I _01706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10459__A1 _04692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09313__A2 _04142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10459__B2 _04514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11120__A2 _04467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07712__B _03132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07875__A2 _03233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11827_ _00523_ net152 u_cpu.rf_ram.memory\[14\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11758_ _00454_ net512 u_cpu.rf_ram.memory\[142\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10709_ u_cpu.rf_ram.memory\[104\]\[2\] _05180_ _05181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11689_ _00393_ net329 u_cpu.rf_ram.memory\[56\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout226_I net228 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11187__A2 _05478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06063__B _01679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06063__A1 _01672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07920_ _03266_ _03255_ _03267_ _00260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09001__A1 _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08769__I _03801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07851_ _03193_ _03216_ _03223_ _00235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10698__A1 _05146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07563__A1 u_cpu.rf_ram.memory\[41\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06610__I0 u_cpu.rf_ram.memory\[96\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06802_ _01740_ _02412_ _02031_ _02413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_111_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06289__I _01675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput2 io_in[1] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07782_ u_cpu.rf_ram.memory\[40\]\[6\] _03172_ _03177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09521_ _03124_ _04286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06733_ u_cpu.rf_ram.memory\[140\]\[5\] u_cpu.rf_ram.memory\[141\]\[5\] u_cpu.rf_ram.memory\[142\]\[5\]
+ u_cpu.rf_ram.memory\[143\]\[5\] _02169_ _01816_ _02345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_77_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11111__A2 _04034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09452_ u_cpu.rf_ram.memory\[115\]\[0\] _04240_ _04241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout41_I net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06664_ _02078_ _02275_ _02276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08403_ _02869_ _03574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11941__CLK net462 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09383_ _02869_ _04198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10870__A1 u_cpu.rf_ram.memory\[108\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06595_ u_cpu.rf_ram.memory\[44\]\[4\] u_cpu.rf_ram.memory\[45\]\[4\] u_cpu.rf_ram.memory\[46\]\[4\]
+ u_cpu.rf_ram.memory\[47\]\[4\] _01692_ _01879_ _02208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_52_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06238__B _01628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08334_ _03498_ _03525_ _03531_ _00410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10475__S _04466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08265_ u_cpu.rf_ram.memory\[57\]\[7\] _03472_ _03483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07216_ _02789_ _02790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08196_ _03438_ _03443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11178__A2 _05477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07147_ u_cpu.cpu.immdec.imm11_7\[4\] _02724_ _02728_ _02729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_88_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09791__A2 _04482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07078_ _02662_ _02660_ _02670_ _00014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05801__A1 _01447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06029_ _01618_ _01629_ _01636_ _01645_ _01428_ _01646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_133_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07554__A1 u_cpu.rf_ram.memory\[41\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12597__CLK net279 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06199__I _01815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09719_ _04437_ _04418_ _04444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_74_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10991_ u_cpu.rf_ram.memory\[110\]\[3\] _05355_ _05358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11102__A2 _01393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[47\]_SE net558 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07857__A2 _03217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12661_ _01340_ net159 u_cpu.rf_ram.memory\[100\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11612_ _00316_ net238 u_cpu.rf_ram.memory\[64\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07959__S _03289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07609__A2 _03052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12592_ _01271_ net278 u_cpu.rf_ram.memory\[88\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11543_ _00247_ net256 u_cpu.rf_ram.memory\[74\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05987__B _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06132__I2 u_cpu.rf_ram.memory\[114\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11474_ _00178_ net110 u_cpu.rf_ram.memory\[4\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06683__I3 u_cpu.rf_ram.memory\[47\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11169__A2 _05466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10184__I _04848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10425_ _04992_ _04994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08034__A2 _03338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10916__A2 _05303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10356_ u_cpu.cpu.ctrl.o_ibus_adr\[30\] _04906_ _04909_ u_cpu.cpu.ctrl.o_ibus_adr\[31\]
+ _04951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_98_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07793__A1 _03179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06596__A2 _02208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11814__CLK net370 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10287_ _04911_ _00984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_26_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06611__B _01663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12026_ _00709_ net490 u_cpu.cpu.state.o_cnt_r\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06348__A2 _01962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07545__A1 _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09922__B _02529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout176_I net184 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07848__A2 _03220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout343_I net344 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06380_ u_cpu.rf_ram.memory\[32\]\[2\] u_cpu.rf_ram.memory\[33\]\[2\] u_cpu.rf_ram.memory\[34\]\[2\]
+ u_cpu.rf_ram.memory\[35\]\[2\] _01705_ _01994_ _01995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout510_I net511 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10455__I1 _02700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08050_ u_cpu.rf_ram.memory\[65\]\[5\] _03343_ _03350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11344__CLK net207 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07001_ u_cpu.cpu.state.o_cnt_r\[2\] u_cpu.cpu.ctrl.i_iscomp _02608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_11_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08025__A2 _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09773__A2 _04485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11494__CLK net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06587__A2 _02199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08952_ _03061_ _03181_ _03921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout89_I net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07903_ u_cpu.rf_ram.memory\[76\]\[0\] _03255_ _03256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08883_ _03874_ _00616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07834_ u_cpu.rf_ram.memory\[129\]\[6\] _03208_ _03213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10391__I0 _04188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09289__A1 u_cpu.rf_ram.memory\[117\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07765_ _03165_ _03166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09504_ u_cpu.rf_ram.memory\[33\]\[2\] _04274_ _04275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06716_ _02147_ _02327_ _02328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07696_ _03117_ _03118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_24_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09435_ _04225_ _04230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10843__A1 _05211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06647_ u_cpu.rf_ram.memory\[128\]\[4\] u_cpu.rf_ram.memory\[129\]\[4\] u_cpu.rf_ram.memory\[130\]\[4\]
+ u_cpu.rf_ram.memory\[131\]\[4\] _01614_ _01827_ _02260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_90_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_94_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_55_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09366_ _04184_ u_cpu.rf_ram.memory\[8\]\[0\] _04186_ _04187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_36_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06578_ _02081_ _02190_ _01970_ _02191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_40_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08317_ u_cpu.rf_ram.memory\[55\]\[5\] _03517_ _03521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09297_ _04141_ _04142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08264__A2 _03474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06275__A1 _01715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10071__A2 _04738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08248_ _03472_ _03473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_125_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06665__I3 u_cpu.rf_ram.memory\[19\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11837__CLK net487 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09213__A1 _03112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08016__A2 _03324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08179_ u_cpu.rf_ram.memory\[60\]\[3\] _03431_ _03433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09793__I _04421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10210_ _04863_ _00955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11020__A1 _05361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11190_ u_cpu.rf_ram.memory\[25\]\[7\] _05476_ _05487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07775__A1 _03071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10141_ _02756_ _04820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09516__A2 _04034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10072_ u_arbiter.i_wb_cpu_rdt\[16\] u_arbiter.i_wb_cpu_rdt\[0\] _01446_ _04760_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10974_ _05284_ _05337_ _05345_ _01237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09033__I _03180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06889__I0 u_cpu.rf_ram.memory\[88\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10834__A1 _05199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06502__A2 _02077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12644_ _01323_ net113 u_cpu.rf_ram.memory\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12612__CLK net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12575_ _01254_ net203 u_cpu.rf_ram.memory\[86\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xu_scanchain_local.scan_flop\[67\] u_scanchain_local.module_data_in\[66\] net554 u_arbiter.o_wb_cpu_adr\[29\]
+ net22 u_scanchain_local.module_data_in\[67\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_8_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08255__A2 _03477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11526_ _00230_ net432 u_cpu.rf_ram.memory\[129\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09204__A1 _01409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08007__A2 _03313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11457_ _00161_ net327 u_cpu.rf_ram.memory\[48\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10408_ _04984_ _01032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11011__A1 _05352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11388_ _00092_ net188 u_cpu.rf_ram.memory\[78\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06569__A2 _02181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06113__S1 _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07766__A1 _03018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10339_ _04941_ _01006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10642__I _05131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout293_I net294 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10117__A3 _04615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12009_ _00692_ net425 u_cpu.rf_ram.memory\[37\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05880_ u_arbiter.i_wb_cpu_dbus_adr\[16\] _01512_ _01513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout460_I net474 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07550_ _03019_ _03020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__11078__A1 _05359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06501_ _01862_ _02102_ _02114_ _02115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_78_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10825__A1 _05213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07481_ _02968_ _02973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08494__A2 _03622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09220_ u_cpu.rf_ram.memory\[92\]\[1\] _04094_ _04096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06432_ _01572_ _02047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_22_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12292__CLK net495 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[43\]_CLK net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09151_ _03969_ _04045_ _04047_ _00711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10817__I _05244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06363_ _01649_ _01977_ _01978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09443__A1 _04154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08246__A2 _03462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08102_ _03381_ _03383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10053__A2 _04636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11250__A1 _02830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09082_ _04002_ _04003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09994__A2 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06294_ _01746_ _01909_ _01910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08033_ _03336_ _03338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08223__S _03450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07757__A1 _03078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10552__I _05083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09984_ u_arbiter.i_wb_cpu_rdt\[27\] u_arbiter.i_wb_cpu_rdt\[11\] _01446_ _04682_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_76_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08935_ _03907_ _03896_ _03908_ _00634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11305__A2 _05548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08866_ _03821_ _03859_ _03864_ _00609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07861__I _03228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08182__A1 _03417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07817_ _03201_ _03202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08797_ _03819_ _03816_ _03820_ _00584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11069__A1 _05347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07748_ _03060_ _03154_ _03156_ _00199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10816__A1 _05204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07679_ _02861_ u_cpu.rf_ram.memory\[4\]\[3\] _03102_ _03106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_41_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09682__A1 _04404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08485__A2 _03625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09788__I _04509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10292__A2 _04907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09418_ _04150_ _04213_ _04219_ _00807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10690_ _05137_ _05164_ _05169_ _01129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09434__A1 _04145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09349_ _04145_ _04173_ _04176_ _00781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08237__A2 _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10044__A2 _04736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12360_ _01039_ net135 u_cpu.rf_ram.memory\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11241__A1 _05454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09985__A2 _04609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07101__I _02690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06638__I3 u_cpu.rf_ram.memory\[79\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11311_ u_cpu.cpu.state.ibus_cyc _05558_ _05559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07996__A1 _03257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12291_ _00022_ net495 u_cpu.cpu.bufreg.c_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11242_ u_cpu.rf_ram.memory\[98\]\[4\] _05515_ _05518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06940__I u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07748__A1 _03060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11173_ _05476_ _05477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10124_ _04804_ _04805_ _04806_ _00926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06420__A1 _01772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12165__CLK net390 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06810__I3 u_cpu.rf_ram.memory\[71\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10055_ u_cpu.cpu.immdec.imm19_12_20\[3\] _04739_ _04745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08173__A1 _03405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07920__A1 _03266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06723__A2 _02334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10957_ _05300_ _02786_ _05335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06487__A1 _02098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10283__A2 _02696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10888_ u_cpu.rf_ram.memory\[69\]\[3\] _05293_ _05295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12627_ _01306_ net54 u_cpu.rf_ram.memory\[25\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09425__A1 u_cpu.rf_ram.memory\[112\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout139_I net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09976__A2 _04672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12558_ _01237_ net212 u_cpu.rf_ram.memory\[85\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06334__S1 _01832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11509_ _00213_ net301 u_cpu.rf_ram.memory\[40\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout306_I net338 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12489_ _01168_ net40 u_cpu.rf_ram.memory\[106\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09728__A2 _04441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07739__A1 _03081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12508__CLK net162 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06981_ u_cpu.cpu.alu.i_rs1 u_cpu.cpu.alu.add_cy_r _02588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06801__I3 u_cpu.rf_ram.memory\[91\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05932_ u_arbiter.i_wb_cpu_dbus_adr\[28\] _01539_ _01553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08720_ u_cpu.rf_ram.memory\[49\]\[4\] _03770_ _03773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11299__A1 _02899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08164__A1 _03421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12658__CLK net160 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08651_ _03676_ _03722_ _03728_ _00530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05863_ u_cpu.cpu.ctrl.o_ibus_adr\[13\] _01495_ _01492_ _01499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_67_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07911__A1 _03259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07602_ _02989_ _03048_ _03053_ _00156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08582_ _03686_ _03687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05794_ _01440_ _01441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_19_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07533_ u_cpu.rf_ram.memory\[51\]\[1\] _03008_ _03010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08467__A2 _03613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11682__CLK net324 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10274__A2 _04898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07464_ _02907_ _02954_ _02961_ _00110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09203_ _04080_ _04082_ _04083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06415_ u_cpu.rf_ram.memory\[88\]\[2\] u_cpu.rf_ram.memory\[89\]\[2\] u_cpu.rf_ram.memory\[90\]\[2\]
+ u_cpu.rf_ram.memory\[91\]\[2\] _02029_ _01768_ _02030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09416__A1 _04147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07395_ _02913_ _02894_ _02914_ _00088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09134_ _04034_ _04035_ _04036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__12038__CLK net285 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10026__A2 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06346_ _01958_ _01960_ _01961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07978__A1 _03259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09065_ _03969_ _03991_ _03993_ _00679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06277_ u_cpu.rf_ram.memory\[104\]\[1\] u_cpu.rf_ram.memory\[105\]\[1\] u_cpu.rf_ram.memory\[106\]\[1\]
+ u_cpu.rf_ram.memory\[107\]\[1\] _01721_ _01892_ _01893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08016_ _03257_ _03324_ _03327_ _00296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09719__A2 _04418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06650__A1 _02060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12188__CLK net390 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10282__I _04906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08888__S _03872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09967_ _04465_ _04666_ _04667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08918_ _02890_ _03814_ _03895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09898_ _04546_ _04453_ _04604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08155__A1 _03415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08849_ u_cpu.rf_ram.memory\[131\]\[4\] _03851_ _03854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06261__S0 _01686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11860_ _00556_ net477 u_cpu.rf_ram.memory\[49\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10811_ _05244_ _05245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11791_ _00487_ net373 u_cpu.rf_ram.memory\[73\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08458__A2 _03610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10265__A2 _04895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10742_ _02922_ _03061_ _05200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09311__I _03909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06859__I3 u_cpu.rf_ram.memory\[47\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10673_ _05142_ _05151_ _05158_ _01123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09407__A1 _02890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07967__S _03288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12412_ _01091_ net81 u_cpu.rf_ram.memory\[28\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09958__A2 _04485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07969__A1 _02831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11405__CLK net221 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10393__S _04973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12343_ _01023_ net165 u_cpu.rf_ram.memory\[109\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12274_ _00957_ net533 u_arbiter.i_wb_cpu_dbus_adr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11225_ _05507_ _01326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11555__CLK net242 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11156_ _05444_ _05465_ _05467_ _01297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_7_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10107_ _04550_ _04791_ _04792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06795__I2 u_cpu.rf_ram.memory\[118\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11087_ _05415_ _05416_ _05417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_27_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10038_ _04608_ _04499_ _04731_ _04585_ _04732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_48_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08697__A2 _03753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09646__A1 u_arbiter.i_wb_cpu_rdt\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout256_I net257 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11989_ _00008_ net263 u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10256__A2 _02705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06200_ u_cpu.rf_ram.memory\[136\]\[0\] u_cpu.rf_ram.memory\[137\]\[0\] u_cpu.rf_ram.memory\[138\]\[0\]
+ u_cpu.rf_ram.memory\[139\]\[0\] _01814_ _01816_ _01817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_13_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11205__A1 _05456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06880__A1 _01672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07180_ u_cpu.rf_ram.memory\[82\]\[3\] _02753_ _02759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06307__S1 _01780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06131_ _01652_ _01748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12330__CLK net504 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08621__A2 _03701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06062_ _01678_ _01679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout406 net407 net406 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_09821_ _04538_ _04539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_99_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12480__CLK net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout417 net424 net417 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_119_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08501__S _03633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout428 net429 net428 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_86_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout439 net440 net439 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05738__A3 _01388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09752_ u_arbiter.i_wb_cpu_rdt\[13\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[13\]
+ _04413_ _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_fanout71_I net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06964_ _02571_ u_cpu.cpu.decode.co_ebreak _01413_ _02572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_100_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08137__A1 _03351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08703_ u_cpu.rf_ram.memory\[137\]\[6\] _03753_ _03762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05915_ u_arbiter.i_wb_cpu_dbus_adr\[24\] _01539_ _01540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08300__I _03509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09683_ _04403_ _04407_ _04408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06895_ _02498_ _02500_ _02502_ _02504_ _01757_ _02505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__08688__A2 _03747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06538__I2 u_cpu.rf_ram.memory\[86\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09840__B _04556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05846_ u_cpu.cpu.ctrl.o_ibus_adr\[9\] _01485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_08634_ _03572_ u_cpu.rf_ram.memory\[14\]\[5\] _03711_ _03718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09637__A1 u_arbiter.i_wb_cpu_rdt\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08565_ _03673_ _03668_ _03675_ _00497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05777_ _01427_ _01428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_35_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout13 net14 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__10247__A2 _02691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07516_ u_cpu.rf_ram.memory\[44\]\[5\] _02990_ _02997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout24 net25 net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08496_ _03632_ _03633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xfanout35 u_scanchain_local.clk net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__06546__S1 _01799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout46 net49 net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_35_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11428__CLK net333 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07447_ u_cpu.rf_ram.memory\[42\]\[6\] _02946_ _02951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout57 net58 net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_10_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout68 net70 net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout79 net83 net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XFILLER_126_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08860__A2 _03860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06871__A1 _01656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07378_ u_cpu.rf_ram.memory\[80\]\[2\] _02901_ _02902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06329_ u_cpu.rf_ram.memory\[140\]\[1\] u_cpu.rf_ram.memory\[141\]\[1\] u_cpu.rf_ram.memory\[142\]\[1\]
+ u_cpu.rf_ram.memory\[143\]\[1\] _01820_ _01821_ _01945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09117_ u_cpu.rf_ram.memory\[36\]\[6\] _04019_ _04024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08612__A2 _03704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06704__B _01679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11578__CLK net349 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09048_ _03980_ _03972_ _03981_ _00674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06423__C _01925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10941__S _05326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11010_ u_cpu.rf_ram.memory\[86\]\[1\] _05369_ _05371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08376__A1 _03501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08411__S _03579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08128__A1 u_cpu.rf_ram.memory\[62\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08210__I _03450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09876__A1 u_cpu.rf_ram.memory\[114\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06529__I2 u_cpu.rf_ram.memory\[94\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06234__S0 _01849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11912_ _00608_ net458 u_cpu.rf_ram.memory\[130\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12203__CLK net384 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11843_ _00539_ net432 u_cpu.rf_ram.memory\[39\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09628__A1 u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11774_ _00470_ net512 u_cpu.rf_ram.memory\[140\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10725_ _05130_ _05188_ _05190_ _01143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12353__CLK net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08851__A2 _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06862__A1 _01715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10656_ _05146_ _05133_ _05147_ _01117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10587_ u_cpu.rf_ram.memory\[28\]\[3\] _05104_ _05106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07496__I _02981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12326_ _01006_ net525 u_cpu.cpu.ctrl.o_ibus_adr\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06465__I1 u_cpu.rf_ram.memory\[21\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12257_ _00940_ net81 u_cpu.rf_ram.memory\[31\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08367__A1 _03485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05945__S _01434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11208_ u_cpu.rf_ram.memory\[24\]\[6\] _05493_ _05498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12188_ _00871_ net390 u_arbiter.i_wb_cpu_dbus_dat\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10174__A1 _04824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06473__S0 _01640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11139_ _05454_ _05446_ _05455_ _01292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08119__A1 _03353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09216__I _04092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07590__A2 _03037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout373_I net374 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10477__A2 _04453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06680_ _02285_ _02287_ _02289_ _02291_ _01427_ _02292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_110_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09619__A1 u_arbiter.i_wb_cpu_rdt\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08350_ _03536_ _03541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09095__A2 _04007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07301_ _02778_ _02834_ _02843_ _00065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08281_ u_cpu.rf_ram.memory\[56\]\[2\] _03495_ _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08842__A2 _03848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07232_ _02768_ _02793_ _02800_ _00039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06853__A1 _01725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07163_ _02735_ u_cpu.rf_ram_if.wdata0_r\[1\] _02743_ _02744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_9_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06605__A1 _02117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06114_ _01662_ _01731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_106_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07094_ _01376_ _02684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06045_ _01601_ _01662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11870__CLK net516 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08358__A1 _03504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout203 net208 net203 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_113_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout214 net230 net214 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__10165__A1 _04808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout225 net228 net225 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_119_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout236 net238 net236 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_09804_ _04436_ _04457_ _04503_ _04521_ _04523_ _04477_ _04524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__07030__A1 u_arbiter.i_wb_cpu_ibus_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout247 net248 net247 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout258 net259 net258 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout269 net540 net269 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__12226__CLK net362 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07996_ _03257_ _03312_ _03315_ _00288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07581__A2 _03040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09735_ _04452_ _04457_ _04459_ _04460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08030__I _03059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06947_ _02553_ _02549_ _02554_ _02555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09858__A1 _02571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06216__S0 _01831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09666_ u_cpu.rf_ram.memory\[113\]\[6\] _04388_ _04393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06878_ _01649_ _02487_ _02488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08530__A1 _03604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08617_ _03680_ _03701_ _03708_ _00516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05829_ u_cpu.cpu.ctrl.o_ibus_adr\[7\] _01468_ _01471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09597_ _04346_ _04348_ _00857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12376__CLK net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06485__I _01675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08548_ _03602_ _03656_ _03663_ _00492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09086__A2 _04004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07097__A1 _02549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08479_ _03588_ _03621_ _03623_ _00463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08833__A2 _03839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09796__I _03118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10510_ _05057_ _05042_ _05058_ _01060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06844__A1 _01590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10640__A2 _05132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11490_ _00194_ net178 u_cpu.rf_ram.memory\[16\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10441_ u_cpu.rf_ram.memory\[93\]\[7\] _04992_ _05003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08597__A1 u_cpu.rf_ram.memory\[70\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10372_ u_cpu.rf_ram.memory\[109\]\[1\] _04962_ _04964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12111_ _00794_ net143 u_cpu.rf_ram.memory\[8\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08349__A1 _03491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09397__I0 _04192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12042_ _00725_ net308 u_cpu.rf_ram.memory\[90\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10156__A1 _04830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09010__A2 _03945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07021__A1 _02569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09849__A1 _04475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08521__A1 u_cpu.rf_ram.memory\[72\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07712__C _02684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11826_ _00522_ net152 u_cpu.rf_ram.memory\[14\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09077__A2 _03995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11743__CLK net256 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11757_ _00453_ net512 u_cpu.rf_ram.memory\[142\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06835__A1 _01580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10708_ _05175_ _05180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11688_ _00392_ net329 u_cpu.rf_ram.memory\[56\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout121_I net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10639_ u_cpu.rf_ram.memory\[101\]\[1\] _05133_ _05136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11893__CLK net468 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout219_I net223 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12309_ _00989_ net523 u_cpu.cpu.ctrl.o_ibus_adr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06694__S0 _02005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout490_I net492 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09001__A2 _03946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10147__A1 u_cpu.rf_ram.memory\[32\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07850_ u_cpu.rf_ram.memory\[139\]\[4\] _03220_ _03223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10698__A2 _05165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06801_ u_cpu.rf_ram.memory\[88\]\[6\] u_cpu.rf_ram.memory\[89\]\[6\] u_cpu.rf_ram.memory\[90\]\[6\]
+ u_cpu.rf_ram.memory\[91\]\[6\] _02029_ _01742_ _02412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_84_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07781_ _03081_ _03169_ _03176_ _00212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput3 io_in[2] net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_09520_ _04284_ _04285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06732_ _01825_ _02343_ _02344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_92_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11111__A3 _04031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09451_ _04238_ _04240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06663_ u_cpu.rf_ram.memory\[20\]\[5\] u_cpu.rf_ram.memory\[21\]\[5\] u_cpu.rf_ram.memory\[22\]\[5\]
+ u_cpu.rf_ram.memory\[23\]\[5\] _01849_ _01965_ _02275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_65_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08402_ _03573_ _00436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09382_ _04197_ _00793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10870__A2 _05276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout34_I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06594_ _01876_ _02206_ _02207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08333_ u_cpu.rf_ram.memory\[54\]\[3\] _03529_ _03531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08815__A2 _03815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08264_ _03421_ _03474_ _03482_ _00389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06826__A1 _02060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07215_ _02701_ _02725_ _02788_ _02789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_08195_ _03410_ _03439_ _03442_ _00360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08579__A1 u_cpu.rf_ram.memory\[71\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07146_ _02727_ _02728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_140_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10386__A1 _04833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09240__A2 _04106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07077_ u_cpu.rf_ram_if.rdata0\[7\] _02665_ _02670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06685__S0 _01716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06028_ _01637_ _01643_ _01644_ _01645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_134_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11616__CLK net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07003__A1 _02564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10689__A2 _05168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07979_ u_cpu.rf_ram.memory\[68\]\[3\] _03303_ _03305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09718_ _04439_ _04442_ _04443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_56_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10990_ _02757_ _05357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11766__CLK net512 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09649_ _04380_ _04322_ _04382_ _00875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_76_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12660_ _01339_ net159 u_cpu.rf_ram.memory\[100\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10861__A2 _05276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11611_ _00315_ net238 u_cpu.rf_ram.memory\[64\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08806__A2 _03822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12591_ _01270_ net206 u_cpu.rf_ram.memory\[87\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11542_ _00246_ net250 u_cpu.rf_ram.memory\[77\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11473_ _00177_ net303 u_cpu.rf_ram.memory\[50\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10424_ _04992_ _04993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09231__A2 _04097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10355_ _04950_ _01013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_83_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10286_ _01431_ _04907_ _04910_ u_arbiter.i_wb_cpu_ibus_adr\[1\] _04911_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[12\] u_arbiter.i_wb_cpu_rdt\[9\] net544 u_arbiter.i_wb_cpu_dbus_dat\[6\]
+ net12 u_arbiter.i_wb_cpu_rdt\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
X_12025_ _00708_ net490 u_cpu.cpu.state.o_cnt_r\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06428__S0 _01792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12541__CLK net293 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08742__A1 u_cpu.rf_ram.memory\[136\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07545__A2 _03008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout169_I net170 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11809_ _00505_ net371 u_cpu.rf_ram.memory\[70\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout503_I net505 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07000_ u_cpu.cpu.state.o_cnt_r\[1\] _02607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_116_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06667__S0 _02084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08981__A1 _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08951_ _03919_ _03897_ _03920_ _00638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07902_ _03253_ _03255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06419__S0 _01773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08882_ _03564_ u_cpu.rf_ram.memory\[12\]\[1\] _03872_ _03874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08733__A1 u_cpu.rf_ram.memory\[136\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07536__A2 _03011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07833_ _03195_ _03205_ _03212_ _00228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10540__A1 _05046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07764_ _02829_ _02936_ _03165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_38_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09503_ _04269_ _04274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06715_ u_cpu.rf_ram.memory\[80\]\[5\] u_cpu.rf_ram.memory\[81\]\[5\] u_cpu.rf_ram.memory\[82\]\[5\]
+ u_cpu.rf_ram.memory\[83\]\[5\] _01651_ _02033_ _02327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07695_ _03115_ u_arbiter.i_wb_cpu_ibus_adr\[1\] _03116_ _03117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_65_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09434_ _04145_ _04226_ _04229_ _00813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06646_ _01819_ _02258_ _01823_ _02259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10843__A2 _05257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_94_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_75_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09365_ _04185_ _04186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_16_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06577_ u_cpu.rf_ram.memory\[16\]\[4\] u_cpu.rf_ram.memory\[17\]\[4\] u_cpu.rf_ram.memory\[18\]\[4\]
+ u_cpu.rf_ram.memory\[19\]\[4\] _01852_ _01968_ _02190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_33_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08316_ _03501_ _03513_ _03520_ _00403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09296_ _03165_ _03970_ _04141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10285__I _04909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08247_ _03380_ _03020_ _03472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[10\]_D u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10359__A1 _04952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08178_ _03412_ _03427_ _03432_ _00353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07129_ _02708_ _02710_ _02711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06658__S0 _01959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11020__A2 _05369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07594__I _03047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10140_ _04817_ _04810_ _04819_ _00929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08972__A1 _02920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07775__A2 _03168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05786__A1 _01431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10071_ _01391_ _04738_ _04758_ _04759_ _00920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_82_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[14\]_SE net542 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08724__A1 u_cpu.rf_ram.memory\[49\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06003__I _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10531__A1 _04091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06938__I _02546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06830__S0 _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09314__I _03912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10973_ u_cpu.rf_ram.memory\[85\]\[6\] _05340_ _05345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10295__B1 _04910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06889__I1 u_cpu.rf_ram.memory\[89\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10834__A2 _05257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06502__A3 _02089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12643_ _01322_ net115 u_cpu.rf_ram.memory\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12094__CLK net408 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12574_ _01253_ net205 u_cpu.rf_ram.memory\[86\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09452__A2 _04240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10195__I _04848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07463__A1 u_cpu.rf_ram.memory\[46\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11525_ _00229_ net430 u_cpu.rf_ram.memory\[129\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[8\]_D u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11456_ _00160_ net370 u_cpu.rf_ram.memory\[48\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09204__A2 _02556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07215__A1 _02701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10407_ _04184_ u_cpu.rf_ram.memory\[2\]\[0\] _04983_ _04984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06649__S0 _02061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11011__A2 _05368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11387_ _00091_ net220 u_cpu.rf_ram.memory\[78\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08963__A1 _03907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07766__A2 _03166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10338_ u_cpu.cpu.ctrl.o_ibus_adr\[22\] _04936_ _04938_ u_cpu.cpu.ctrl.o_ibus_adr\[23\]
+ _04941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10269_ _04817_ _04894_ _04899_ _00978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07009__I _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09912__B1 _04561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12008_ _00691_ net409 u_cpu.rf_ram.memory\[37\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10522__A1 _05049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout286_I net288 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06821__S0 _02169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout453_I net455 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10286__B1 _04910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06500_ _02105_ _02108_ _02111_ _02113_ _01711_ _02114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_46_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07480_ _02897_ _02969_ _02972_ _00115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10825__A2 _05246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12437__CLK net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06431_ _01797_ _02045_ _02046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09150_ u_cpu.rf_ram.memory\[91\]\[0\] _04046_ _04047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06362_ u_cpu.rf_ram.memory\[52\]\[2\] u_cpu.rf_ram.memory\[53\]\[2\] u_cpu.rf_ram.memory\[54\]\[2\]
+ u_cpu.rf_ram.memory\[55\]\[2\] _01863_ _01653_ _01977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_33_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10589__A1 u_cpu.rf_ram.memory\[28\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09443__A2 _04227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08101_ _03381_ _03382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12587__CLK net200 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06293_ u_cpu.rf_ram.memory\[112\]\[1\] u_cpu.rf_ram.memory\[113\]\[1\] u_cpu.rf_ram.memory\[114\]\[1\]
+ u_cpu.rf_ram.memory\[115\]\[1\] _01747_ _01908_ _01909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__11250__A2 _04958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09081_ _02785_ _02940_ _04002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08032_ _03336_ _03337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_122_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09827__C _04486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[37\]_SE net556 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07757__A2 _03154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09983_ _04468_ _04566_ _04523_ _04680_ _04486_ _04681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_89_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08934_ u_cpu.rf_ram.memory\[128\]\[3\] _03904_ _03908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06280__I2 u_cpu.rf_ram.memory\[102\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08706__A1 u_cpu.rf_ram.memory\[137\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06980__A3 _02586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08865_ u_cpu.rf_ram.memory\[130\]\[2\] _03863_ _03864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07816_ _02724_ _02727_ _03201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_79_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12700__D u_cpu.rf_ram_if.wdata1_r\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06812__S0 _01762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08796_ u_cpu.rf_ram.memory\[133\]\[1\] _03817_ _03820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07747_ u_cpu.rf_ram.memory\[17\]\[0\] _03155_ _03156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05940__A1 u_arbiter.i_wb_cpu_dbus_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09131__A1 _04031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08973__I _03933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10816__A2 _05245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07678_ _03105_ _00180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09682__A2 u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09417_ u_cpu.rf_ram.memory\[112\]\[3\] _04217_ _04219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06629_ u_cpu.rf_ram.memory\[84\]\[4\] u_cpu.rf_ram.memory\[85\]\[4\] u_cpu.rf_ram.memory\[86\]\[4\]
+ u_cpu.rf_ram.memory\[87\]\[4\] _01922_ _02151_ _02242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_41_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09348_ u_cpu.rf_ram.memory\[121\]\[1\] _04174_ _04176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06493__I _01417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09434__A2 _04226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06879__S0 _01674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07445__A1 u_cpu.rf_ram.memory\[42\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09279_ _04056_ _04129_ _04131_ _00756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11241__A2 _05511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11310_ _04511_ _04037_ _05558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07996__A2 _03312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12290_ _00973_ net501 u_arbiter.i_wb_cpu_dbus_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11954__CLK net440 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11241_ _05454_ _05511_ _05517_ _01332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06442__B _01823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07748__A2 _03154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11172_ _05098_ _03020_ _05476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10752__A1 u_cpu.rf_ram.memory\[79\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10123_ u_cpu.cpu.genblk3.csr.mie_mtie u_cpu.cpu.genblk3.csr.mstatus_mie u_cpu.cpu.genblk3.csr.i_mtip
+ _04805_ _04806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__06420__A2 _02034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10054_ _04743_ _04738_ _04744_ _04537_ _00918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_23_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10504__A1 _05053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[5\] u_arbiter.i_wb_cpu_rdt\[2\] net548 u_arbiter.i_wb_cpu_dbus_sel\[3\]
+ net15 u_arbiter.i_wb_cpu_rdt\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_87_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06803__S0 _01651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07920__A2 _03255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09122__A1 _04026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10807__A2 _05231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10956_ _05334_ _01230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11484__CLK net378 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06731__I0 u_cpu.rf_ram.memory\[136\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10887_ _05275_ _05289_ _05294_ _01201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_43_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12626_ _01305_ net53 u_cpu.rf_ram.memory\[25\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12557_ _01236_ net212 u_cpu.rf_ram.memory\[85\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07987__A2 _03298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11508_ _00212_ net303 u_cpu.rf_ram.memory\[40\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12488_ _01167_ net41 u_cpu.rf_ram.memory\[106\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout201_I net202 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11439_ _00143_ net330 u_cpu.rf_ram.memory\[41\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05747__I _01397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07739__A2 _03143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09984__I0 u_arbiter.i_wb_cpu_rdt\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06980_ _02553_ _02585_ _02586_ _02587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05931_ u_cpu.cpu.ctrl.o_ibus_adr\[28\] _01551_ _01552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11299__A2 _05547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08164__A2 _03408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08650_ u_cpu.rf_ram.memory\[138\]\[3\] _03726_ _03728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05862_ _01495_ _01492_ u_cpu.cpu.ctrl.o_ibus_adr\[13\] _01498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_113_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07911__A2 _03254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07601_ u_cpu.rf_ram.memory\[48\]\[2\] _03052_ _03053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08581_ _03272_ _03287_ _03686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05793_ _01439_ _01440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11827__CLK net152 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09113__A1 u_cpu.rf_ram.memory\[36\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07532_ _02980_ _03007_ _03009_ _00130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09664__A2 _04388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07463_ u_cpu.rf_ram.memory\[46\]\[4\] _02958_ _02961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09202_ _02551_ _04081_ _04082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06414_ _01704_ _02029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_50_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11977__CLK net265 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07394_ u_cpu.rf_ram.memory\[80\]\[6\] _02901_ _02914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07202__I _02776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09133_ _04031_ _04030_ _04035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06345_ u_cpu.rf_ram.memory\[4\]\[2\] u_cpu.rf_ram.memory\[5\]\[2\] u_cpu.rf_ram.memory\[6\]\[2\]
+ u_cpu.rf_ram.memory\[7\]\[2\] _01959_ _01592_ _01960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_124_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07978__A2 _03299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09064_ u_cpu.rf_ram.memory\[38\]\[0\] _03992_ _03993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06276_ _01659_ _01892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10982__A1 _05347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08015_ u_cpu.rf_ram.memory\[66\]\[1\] _03325_ _03327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06650__A2 _02262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09129__I _01432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10734__A1 _05142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06402__A2 _02016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09966_ _02529_ _04665_ _04666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06253__I2 u_cpu.rf_ram.memory\[62\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11357__CLK net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12602__CLK net373 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08917_ _03893_ _03894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09897_ _04403_ _04602_ _04603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09352__A1 _04147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08155__A2 _03407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08848_ _03824_ _03847_ _03853_ _00602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06166__A1 _01778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05913__A1 _01537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08779_ _03755_ _03802_ _03808_ _00578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06261__S1 _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09104__A1 u_cpu.rf_ram.memory\[36\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10810_ _03033_ _05243_ _05244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11790_ _00486_ net347 u_cpu.rf_ram.memory\[72\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09655__A2 _04385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07313__S _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10741_ _04807_ _05199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06469__A2 _02082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07666__A1 _03081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06713__I0 u_cpu.rf_ram.memory\[88\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10672_ u_cpu.rf_ram.memory\[102\]\[4\] _05155_ _05158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07112__I _02674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09407__A2 _03970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12411_ _01090_ net90 u_cpu.rf_ram.memory\[28\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07969__A2 _02923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06951__I _01371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12342_ _01022_ net165 u_cpu.rf_ram.memory\[109\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08091__A1 u_cpu.rf_ram.memory\[29\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12132__CLK net436 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12273_ _00956_ net531 u_arbiter.i_wb_cpu_dbus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06641__A2 _02244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09039__I _03899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08918__A1 _02890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11224_ _02866_ u_cpu.rf_ram.memory\[0\]\[5\] _05500_ _05507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10725__A1 _05130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11155_ u_cpu.rf_ram.memory\[26\]\[0\] _05466_ _05467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12282__CLK net525 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10106_ _04650_ _04710_ _04791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06795__I3 u_cpu.rf_ram.memory\[119\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11086_ _02529_ _02572_ _02565_ _05416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_27_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09343__A1 _03019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10037_ _04729_ _04730_ _04731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_76_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11150__A1 u_cpu.rf_ram.memory\[27\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09894__A2 _04599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[57\]_CLK net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11988_ _00678_ net439 u_cpu.rf_ram.memory\[123\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07657__A1 _03068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout151_I net155 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10939_ _03870_ _02938_ _05325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_56_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout249_I net255 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12609_ _01288_ net380 u_cpu.cpu.genblk3.csr.o_new_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07409__A1 u_cpu.rf_ram.memory\[78\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06880__A2 _02489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout416_I net417 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06130_ _01650_ _01747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_118_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08082__A1 u_cpu.rf_ram.memory\[29\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06061_ _01417_ _01678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08909__A1 _03826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10716__A1 _05144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09820_ _04421_ _04423_ _04506_ _04538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_99_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout407 net413 net407 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_98_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout418 net424 net418 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__08788__I _03484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout429 net433 net429 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_101_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09751_ _04431_ _04475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_45_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06963_ u_cpu.cpu.decode.op21 _02571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_67_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08702_ _03506_ _03761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09334__A1 _04150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08137__A2 _03395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05914_ _01451_ _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09682_ _04404_ u_arbiter.i_wb_cpu_rdt\[8\] _04406_ _04407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_80_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06148__A1 _01761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout64_I net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06894_ _02150_ _02503_ _02153_ _02504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11141__A1 u_cpu.rf_ram.memory\[27\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08633_ _03717_ _00523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05845_ u_cpu.cpu.ctrl.o_ibus_adr\[10\] _01484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07896__A1 _03197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06699__A2 _02310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08564_ u_cpu.rf_ram.memory\[71\]\[2\] _03674_ _03675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12005__CLK net408 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05776_ _01426_ _01427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09637__A2 _04293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07515_ _02909_ _02996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_93_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10558__I _05083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout14 net19 net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_08495_ _03285_ _02967_ _03632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_126_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout25 net33 net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_39_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout36 u_arbiter.i_wb_cpu_dbus_dat\[1\] net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout47 net48 net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_126_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07446_ _02910_ _02943_ _02950_ _00103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout58 net61 net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_91_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout69 net70 net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_10_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06871__A2 _02480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07377_ _02892_ _02901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09116_ _03984_ _04016_ _04023_ _00700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08073__A1 _03349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06328_ _01400_ _01943_ _01944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_87_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09047_ u_cpu.rf_ram.memory\[123\]\[3\] _03978_ _03981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06259_ _01865_ _01868_ _01870_ _01874_ _01681_ _01875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_85_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10707__A1 _05135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08376__A2 _03549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09949_ _04504_ _04650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_63_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11132__A1 _05449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11911_ _00607_ net457 u_cpu.rf_ram.memory\[130\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06011__I _01627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06234__S1 _01616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11842_ _00538_ net432 u_cpu.rf_ram.memory\[39\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09628__A2 _04295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11773_ _00469_ net514 u_cpu.rf_ram.memory\[140\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07103__A3 _02635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10724_ u_cpu.rf_ram.memory\[99\]\[0\] _05189_ _05190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10655_ u_cpu.rf_ram.memory\[101\]\[6\] _05138_ _05147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06862__A2 _02471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08064__A1 _03340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11522__CLK net430 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12648__CLK net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10586_ _05046_ _05100_ _05105_ _01089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_12325_ _01005_ net526 u_cpu.cpu.ctrl.o_ibus_adr\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xu_scanchain_local.scan_flop\[42\] u_scanchain_local.module_data_in\[41\] net553 u_arbiter.o_wb_cpu_adr\[4\]
+ net21 u_scanchain_local.module_data_in\[42\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_86_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07811__A1 u_cpu.rf_ram.memory\[119\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06614__A2 _02226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06465__I2 u_cpu.rf_ram.memory\[22\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12256_ _00939_ net93 u_cpu.rf_ram.memory\[31\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09564__A1 u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11672__CLK net314 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08367__A2 _03549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11207_ _05458_ _05490_ _05497_ _01318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_12187_ _00870_ net497 u_arbiter.i_wb_cpu_dbus_dat\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10174__A2 _04836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11138_ u_cpu.rf_ram.memory\[27\]\[3\] _05452_ _05455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06473__S1 _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09316__A1 _04154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08119__A2 _03383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12028__CLK net320 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11069_ _05347_ _05404_ _05406_ _01271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11123__A1 _03111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07878__A1 _03199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout366_I net367 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09619__A2 _04311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12178__CLK net386 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout533_I net534 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07300_ u_cpu.rf_ram.memory\[20\]\[7\] _02832_ _02843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08280_ _03486_ _03495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07350__I0 _02858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07231_ u_cpu.rf_ram.memory\[21\]\[5\] _02796_ _02800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10237__I0 u_arbiter.i_wb_cpu_dbus_adr\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07162_ _02736_ u_cpu.rf_ram_if.wdata1_r\[1\] _02743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_30_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10937__A1 u_cpu.rf_ram.memory\[59\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06113_ u_cpu.rf_ram.memory\[96\]\[0\] u_cpu.rf_ram.memory\[97\]\[0\] u_cpu.rf_ram.memory\[98\]\[0\]
+ u_cpu.rf_ram.memory\[99\]\[0\] _01729_ _01641_ _01730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07093_ _02549_ u_cpu.cpu.bufreg.c_r _02681_ _02682_ _02683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_12_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07802__A1 u_cpu.rf_ram.memory\[119\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11002__I _02777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06044_ u_cpu.rf_ram.memory\[48\]\[0\] u_cpu.rf_ram.memory\[49\]\[0\] u_cpu.rf_ram.memory\[50\]\[0\]
+ u_cpu.rf_ram.memory\[51\]\[0\] _01657_ _01660_ _01661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_86_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08358__A2 _03538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout204 net208 net204 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_82_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06369__A1 _01672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout215 net219 net215 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_86_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10165__A2 _04836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout226 net228 net226 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_09803_ _04522_ _04523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout237 net238 net237 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_8_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07030__A2 _02635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout248 net267 net248 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__10062__B _04750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07995_ u_cpu.rf_ram.memory\[67\]\[1\] _03313_ _03315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout259 net260 net259 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_75_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09307__A1 _04147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09734_ _04458_ _04459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06946_ _02553_ _01391_ _02554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09858__A2 _04398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09665_ _04251_ _04385_ _04392_ _00881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06216__S1 _01832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06877_ u_cpu.rf_ram.memory\[124\]\[7\] u_cpu.rf_ram.memory\[125\]\[7\] u_cpu.rf_ram.memory\[126\]\[7\]
+ u_cpu.rf_ram.memory\[127\]\[7\] _01773_ _01774_ _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_27_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08530__A2 _03644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08616_ u_cpu.rf_ram.memory\[143\]\[5\] _03704_ _03708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05828_ _01467_ _01469_ _01470_ u_arbiter.o_wb_cpu_adr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_93_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09596_ u_arbiter.i_wb_cpu_rdt\[13\] _04347_ _04344_ u_arbiter.i_wb_cpu_dbus_dat\[13\]
+ _04348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08547_ u_cpu.rf_ram.memory\[73\]\[5\] _03659_ _03663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05759_ u_cpu.cpu.decode.co_mem_word u_cpu.cpu.bne_or_bge _01410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_70_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11545__CLK net258 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08294__A1 _03504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08478_ u_cpu.rf_ram.memory\[140\]\[0\] _03622_ _03623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07429_ _02700_ _02788_ _02847_ _02939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_17_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06844__A2 _02453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10440_ _04830_ _04994_ _05002_ _01046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10928__A1 _05275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09794__A1 _02676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08597__A2 _03691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10371_ _04808_ _04961_ _04963_ _01016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06152__S0 _01767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12110_ _00793_ net127 u_cpu.rf_ram.memory\[8\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06006__I u_cpu.raddr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09546__A1 u_arbiter.i_wb_cpu_rdt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08349__A2 _03537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12041_ _00724_ net308 u_cpu.rf_ram.memory\[90\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10156__A2 _04811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09317__I _03915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07021__A2 _02625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11105__A1 _04026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09849__A2 _04490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10399__S _04972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06907__I0 u_cpu.rf_ram.memory\[136\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12320__CLK net532 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08521__A2 _03647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06532__A1 _01766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09052__I _03912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11825_ _00521_ net149 u_cpu.rf_ram.memory\[14\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11756_ _00452_ net512 u_cpu.rf_ram.memory\[142\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08285__A1 u_cpu.rf_ram.memory\[56\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10092__A1 _04692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10707_ _05135_ _05176_ _05179_ _01136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06835__A2 _02444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11687_ _00391_ net329 u_cpu.rf_ram.memory\[56\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06391__S0 _02005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10638_ _04813_ _05135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_127_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10919__A1 _03004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09785__A1 _04503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout114_I net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10569_ u_cpu.rf_ram.memory\[96\]\[7\] _05083_ _05094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12308_ _00988_ net523 u_cpu.cpu.ctrl.o_ibus_adr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06694__S1 _01892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12239_ _00922_ net341 u_cpu.cpu.immdec.imm19_12_20\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10661__I _05150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout483_I net484 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11418__CLK net291 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06800_ _01735_ _02410_ _02411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08760__A2 _03794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06610__I2 u_cpu.rf_ram.memory\[98\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07780_ u_cpu.rf_ram.memory\[40\]\[5\] _03172_ _03176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07970__I _03298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput4 io_in[3] net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_37_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06731_ u_cpu.rf_ram.memory\[136\]\[5\] u_cpu.rf_ram.memory\[137\]\[5\] u_cpu.rf_ram.memory\[138\]\[5\]
+ u_cpu.rf_ram.memory\[139\]\[5\] _01831_ _01942_ _02343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_42_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11111__A4 _02562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09450_ _04238_ _04239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_92_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06662_ _02267_ _02269_ _02271_ _02273_ _01807_ _02274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11568__CLK net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08401_ _03572_ u_cpu.rf_ram.memory\[9\]\[5\] _03561_ _03573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_24_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09381_ _04196_ u_cpu.rf_ram.memory\[8\]\[5\] _04185_ _04197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_17_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06593_ u_cpu.rf_ram.memory\[40\]\[4\] u_cpu.rf_ram.memory\[41\]\[4\] u_cpu.rf_ram.memory\[42\]\[4\]
+ u_cpu.rf_ram.memory\[43\]\[4\] _01686_ _02103_ _02206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_52_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08332_ _03494_ _03525_ _03530_ _00409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08276__A1 u_cpu.rf_ram.memory\[56\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout27_I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08507__S _03632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07323__I0 _02861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08263_ u_cpu.rf_ram.memory\[57\]\[6\] _03477_ _03482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06826__A2 _02436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07214_ _02787_ _02728_ _02788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_14_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08194_ u_cpu.rf_ram.memory\[19\]\[1\] _03440_ _03442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07145_ _02726_ u_cpu.rf_ram_if.wen1_r u_cpu.rf_ram_if.rtrig0 u_cpu.rf_ram_if.wen0_r
+ _02727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_106_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10386__A2 _04962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10630__I0 u_arbiter.i_wb_cpu_rdt\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07076_ _02662_ _02658_ _02669_ _00013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07251__A2 _02810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06685__S1 _02109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12703__D u_cpu.rf_ram_if.wdata1_r\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06027_ _01418_ _01644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06270__B _01709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08200__A1 _03415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08751__A2 _03791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07978_ _03259_ _03299_ _03304_ _00281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_59_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09717_ _04441_ _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06929_ u_arbiter.i_wb_cpu_dbus_we _02536_ u_cpu.cpu.immdec.imm24_20\[0\] _02538_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_74_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09648_ u_arbiter.i_wb_cpu_rdt\[31\] _04290_ _04371_ _02547_ _04382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_95_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06514__A1 _02119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09579_ _04333_ _04335_ _00852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10947__S _05326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11610_ _00314_ net237 u_cpu.rf_ram.memory\[64\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12590_ _01269_ net206 u_cpu.rf_ram.memory\[87\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08417__S _03579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07321__S _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10074__A1 _04602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11541_ _00245_ net249 u_cpu.rf_ram.memory\[77\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06817__A2 _02418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08019__A1 _03259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11472_ _00176_ net346 u_cpu.rf_ram.memory\[50\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07490__A2 _02973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10423_ _04091_ _02967_ _04992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09756__B _04479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10377__A2 _04965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10354_ u_cpu.cpu.ctrl.o_ibus_adr\[29\] _04906_ _04945_ u_cpu.cpu.ctrl.o_ibus_adr\[30\]
+ _04950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07242__A2 _02807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06676__S1 _01633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08990__A2 _03933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10285_ _04909_ _04910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_3_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12024_ _00707_ net482 u_cpu.cpu.state.o_cnt_r\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06428__S1 _01930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08742__A2 _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11710__CLK net416 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06505__A1 _02117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11860__CLK net477 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11808_ _00504_ net376 u_cpu.rf_ram.memory\[70\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08258__A1 _03415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10065__A1 _04601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11739_ _00443_ net152 u_cpu.rf_ram.memory\[15\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout231_I net268 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout329_I net332 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06364__S0 _01657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07233__A2 _02796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06667__S1 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12366__CLK net210 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08981__A2 _03934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08950_ u_cpu.rf_ram.memory\[128\]\[7\] _03895_ _03920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11317__A1 _04032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06992__A1 u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07901_ _03253_ _03254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08881_ _03873_ _00615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06419__S1 _02033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07832_ u_cpu.rf_ram.memory\[129\]\[5\] _03208_ _03212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09930__B2 u_cpu.cpu.immdec.imm24_20\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10540__A2 _05072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11390__CLK net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07763_ _03087_ _03155_ _03164_ _00206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09502_ _04242_ _04270_ _04273_ _00837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06714_ _01740_ _02325_ _02031_ _02326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07694_ net8 _01433_ _03116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_65_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09433_ u_cpu.rf_ram.memory\[122\]\[1\] _04227_ _04229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06645_ u_cpu.rf_ram.memory\[140\]\[4\] u_cpu.rf_ram.memory\[141\]\[4\] u_cpu.rf_ram.memory\[142\]\[4\]
+ u_cpu.rf_ram.memory\[143\]\[4\] _02169_ _01816_ _02258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_94_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06898__I2 u_cpu.rf_ram.memory\[70\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_94_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09364_ _03870_ _03166_ _04185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_24_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06576_ _02078_ _02188_ _02189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10056__A1 u_cpu.cpu.csr_imm vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08315_ u_cpu.rf_ram.memory\[55\]\[4\] _03517_ _03520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09997__A1 _04494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09295_ _03893_ _04140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06265__B _01695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08246_ _03423_ _03462_ _03471_ _00382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08036__I _03067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07472__A2 _02919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06680__B1 _02289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08177_ u_cpu.rf_ram.memory\[60\]\[2\] _03431_ _03432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07128_ _02535_ _02709_ _02710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06658__S1 _02071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07059_ _02647_ _02658_ _02659_ _00019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08972__A2 _03181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06983__A1 _01412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05786__A2 _01434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11733__CLK net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10070_ u_cpu.cpu.immdec.imm19_12_20\[5\] _04630_ _04739_ _04759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10531__A2 _03062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06586__I1 u_cpu.rf_ram.memory\[49\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06830__S1 _01592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08488__A1 _03600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10972_ _05282_ _05337_ _05344_ _01236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10295__B2 _01463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12642_ _01321_ net112 u_cpu.rf_ram.memory\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12239__CLK net341 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09330__I _04160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09988__A1 _04684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12573_ _01252_ net205 u_cpu.rf_ram.memory\[86\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11524_ _00228_ net432 u_cpu.rf_ram.memory\[129\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08660__A1 _02876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12389__CLK net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11455_ _00159_ net370 u_cpu.rf_ram.memory\[48\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06903__B _01770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10406_ _04982_ _04983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06649__S1 _02174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11386_ _00090_ net220 u_cpu.rf_ram.memory\[78\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10337_ _04940_ _01005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08963__A2 _03922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06974__A1 u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10268_ u_cpu.rf_ram.memory\[30\]\[2\] _04898_ _04899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09912__A1 _04608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12007_ _00690_ net409 u_cpu.rf_ram.memory\[37\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09912__B2 _04601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10199_ _04857_ _00950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10522__A2 _05060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout181_I net183 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06821__S1 _01816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout279_I net280 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08479__A1 _03588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10286__A1 _01431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10286__B2 u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout446_I net447 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06430_ u_cpu.rf_ram.memory\[72\]\[2\] u_cpu.rf_ram.memory\[73\]\[2\] u_cpu.rf_ram.memory\[74\]\[2\]
+ u_cpu.rf_ram.memory\[75\]\[2\] _01934_ _01799_ _02045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_62_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10038__A1 _04608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10038__B2 _04585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09979__A1 _04425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06361_ _01967_ _01971_ _01973_ _01975_ _01428_ _01976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__11606__CLK net244 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10589__A2 _05104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08100_ _03380_ _03062_ _03381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09080_ _03988_ _03992_ _04001_ _00686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08651__A1 _03676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06292_ _01652_ _01908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08031_ _02804_ _02923_ _03336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11756__CLK net512 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09982_ _04602_ _04680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout94_I net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06965__A1 _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10761__A2 _05207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08933_ _03906_ _03907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06104__I _01620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09903__A1 _04489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08864_ _03858_ _03863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07815_ _03199_ _03184_ _03200_ _00222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10070__B _04739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06812__S1 _01763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08795_ _03490_ _03819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07746_ _03153_ _03155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05940__A2 _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10277__A1 _04830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07677_ _02858_ u_cpu.rf_ram.memory\[4\]\[2\] _03102_ _03105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_26_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09416_ _04147_ _04213_ _04218_ _00806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06628_ _02147_ _02240_ _02241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09347_ _04140_ _04173_ _04175_ _00780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06559_ _01947_ _02172_ _02173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12531__CLK net271 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09278_ u_cpu.rf_ram.memory\[117\]\[0\] _04130_ _04131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07445__A2 _02946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06879__S1 _01676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08229_ _03460_ _03462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11240_ u_cpu.rf_ram.memory\[98\]\[3\] _05515_ _05517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12681__CLK net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06256__I0 u_cpu.rf_ram.memory\[56\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11171_ _05462_ _05466_ _05475_ _01304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10752__A2 _05207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10122_ _04026_ _02705_ _04805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__06014__I _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10053_ u_cpu.cpu.immdec.imm19_12_20\[3\] _04636_ _04737_ _04744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_114_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06949__I _01372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06708__A1 _01691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09325__I _04160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10504__A2 _05042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06803__S1 _02033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09122__A2 _03123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10955_ _04200_ u_cpu.rf_ram.memory\[10\]\[7\] _05325_ _05334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07133__A1 _02578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10200__S _04855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10886_ u_cpu.rf_ram.memory\[69\]\[2\] _05293_ _05294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06731__I1 u_cpu.rf_ram.memory\[137\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12625_ _01304_ net57 u_cpu.rf_ram.memory\[26\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06319__S0 _01934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12556_ _01235_ net213 u_cpu.rf_ram.memory\[85\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09928__C _04557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10440__A1 _04830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11507_ _00211_ net302 u_cpu.rf_ram.memory\[40\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12487_ _01166_ net48 u_cpu.rf_ram.memory\[105\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11438_ _00142_ net330 u_cpu.rf_ram.memory\[41\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09984__I1 u_arbiter.i_wb_cpu_rdt\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11369_ _00073_ net133 u_cpu.rf_ram.memory\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06947__A1 _02553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05930_ _01547_ _01548_ _01551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12404__CLK net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05861_ _01473_ _01496_ _01497_ u_arbiter.o_wb_cpu_adr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout563_I net564 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07600_ _03047_ _03052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08580_ _03684_ _03669_ _03685_ _00502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05792_ _01438_ _01439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_82_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09113__A2 _04019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07531_ u_cpu.rf_ram.memory\[51\]\[0\] _03008_ _03009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06558__S0 _01826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12554__CLK net212 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07462_ _02904_ _02954_ _02960_ _00109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_90_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08872__A1 _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09201_ _02547_ _04079_ _04081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_91_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06413_ _01761_ _02027_ _02028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07393_ _02912_ _02913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09132_ u_cpu.cpu.mem_bytecnt\[1\] _04034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06344_ _01787_ _01959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__07427__A2 _02936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06486__I0 u_cpu.rf_ram.memory\[56\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09063_ _03990_ _03992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06275_ _01715_ _01890_ _01891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08014_ _03252_ _03324_ _03326_ _00295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10982__A2 _05349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06789__I1 u_cpu.rf_ram.memory\[125\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09965_ _02679_ _02703_ _02677_ _04665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_98_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08916_ _02738_ _03893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09896_ _04454_ _04602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10498__A1 _05049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09352__A2 _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08847_ u_cpu.rf_ram.memory\[131\]\[3\] _03851_ _03853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[11\]_SI u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08778_ u_cpu.rf_ram.memory\[134\]\[3\] _03806_ _03808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05913__A2 _01535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07729_ u_cpu.rf_ram.memory\[16\]\[1\] _03143_ _03145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10740_ _05148_ _05189_ _05198_ _01150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_41_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08863__A1 _03819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06713__I1 u_cpu.rf_ram.memory\[89\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10670__A1 u_cpu.rf_ram.memory\[102\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10955__S _05325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10671_ _05140_ _05151_ _05157_ _01122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_41_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12410_ _01089_ net90 u_cpu.rf_ram.memory\[28\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08615__A1 _03678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07418__A2 _02929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08425__S _03578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12341_ _01021_ net165 u_cpu.rf_ram.memory\[109\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10973__A2 _05340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12272_ _00955_ net531 u_arbiter.i_wb_cpu_dbus_adr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11222__I0 _02863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11223_ _05506_ _01325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08918__A2 _03814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09040__A1 u_cpu.rf_ram.memory\[123\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06929__A1 u_arbiter.i_wb_cpu_dbus_we vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11154_ _05464_ _05466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_49_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10105_ _04772_ _04788_ _04789_ _04790_ _00923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_62_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11085_ _04026_ _02579_ _05415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09055__I _03915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10036_ _04436_ _04510_ _04652_ _04608_ _04582_ _04730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_76_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09343__A2 _03970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12577__CLK net168 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11451__CLK net333 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11150__A2 _05445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11987_ _00677_ net439 u_cpu.rf_ram.memory\[123\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[27\]_SE net547 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10938_ _05286_ _05315_ _05324_ _01222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08854__A1 _03830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07657__A2 _03090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout144_I net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10869_ _04826_ _05282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_73_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12608_ _01287_ net360 u_cpu.cpu.ctrl.i_iscomp vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08606__A1 _03666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07409__A2 _02926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout311_I net315 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12539_ _01218_ net293 u_cpu.rf_ram.memory\[59\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08082__A2 _03370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_fanout409_I net412 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05758__I _01408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06093__A1 _01703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06060_ u_cpu.rf_ram.memory\[56\]\[0\] u_cpu.rf_ram.memory\[57\]\[0\] u_cpu.rf_ram.memory\[58\]\[0\]
+ u_cpu.rf_ram.memory\[59\]\[0\] _01674_ _01676_ _01677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_99_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08909__A2 _03882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09031__A1 _03919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10716__A2 _05177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout408 net412 net408 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout419 net423 net419 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA_u_scanchain_local.scan_flop\[34\]_SI u_arbiter.i_wb_cpu_dbus_dat\[28\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07593__A1 _02891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09750_ _04473_ _04474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06962_ _02569_ u_cpu.cpu.genblk3.csr.mcause31 _02564_ _02570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_140_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05913_ _01537_ _01535_ _01538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08701_ _03759_ _03748_ _03760_ _00548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09334__A2 _04161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09681_ _04405_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[8\] _04406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06893_ u_cpu.rf_ram.memory\[84\]\[7\] u_cpu.rf_ram.memory\[85\]\[7\] u_cpu.rf_ram.memory\[86\]\[7\]
+ u_cpu.rf_ram.memory\[87\]\[7\] _01752_ _02151_ _02503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_95_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11141__A2 _05452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08632_ _03570_ u_cpu.rf_ram.memory\[14\]\[4\] _03712_ _03717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05844_ u_arbiter.i_wb_cpu_dbus_adr\[10\] _01453_ _01483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07896__A2 _03242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout57_I net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11944__CLK net461 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08563_ _03667_ _03674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05775_ _01424_ _01425_ _01426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_81_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09098__A1 _03986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07514_ _02994_ _02984_ _02995_ _00126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_93_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08494_ _03606_ _03622_ _03631_ _00470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09893__I0 u_arbiter.i_wb_cpu_rdt\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout15 net16 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout26 net28 net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07213__I u_cpu.cpu.immdec.imm11_7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout37 net43 net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__06856__B1 _02463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07445_ u_cpu.rf_ram.memory\[42\]\[5\] _02946_ _02950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout48 net49 net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_23_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout59 net61 net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_126_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06320__A2 _01935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07376_ _02899_ _02900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09115_ u_cpu.rf_ram.memory\[36\]\[5\] _04019_ _04023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06327_ u_cpu.rf_ram.memory\[136\]\[1\] u_cpu.rf_ram.memory\[137\]\[1\] u_cpu.rf_ram.memory\[138\]\[1\]
+ u_cpu.rf_ram.memory\[139\]\[1\] _01814_ _01942_ _01943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_17_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09270__A1 _04070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06703__S0 _01674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06273__B _01888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09046_ _03906_ _03980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06258_ _01672_ _01872_ _01873_ _01874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_136_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05831__A1 _01456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06189_ _01802_ _01804_ _01805_ _01806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08979__I _03933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10707__A2 _05176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07959__I0 _02861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11474__CLK net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07584__A1 _02992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09948_ _04629_ _04647_ _04648_ _04649_ _00907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_24_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09879_ _04242_ _04588_ _04591_ _00896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11910_ _00606_ net457 u_cpu.rf_ram.memory\[131\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10340__B1 _04938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07887__A2 _03245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09603__I _04318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10891__A1 _05280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09089__A1 u_cpu.rf_ram.memory\[37\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11841_ _00537_ net422 u_cpu.rf_ram.memory\[39\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06448__B _01419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11772_ _00468_ net514 u_cpu.rf_ram.memory\[140\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08836__A1 _03832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10723_ _05187_ _05189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06698__I0 u_cpu.rf_ram.memory\[96\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10654_ _04829_ _05146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_70_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08064__A2 _03356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09261__A1 _04061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10585_ u_cpu.rf_ram.memory\[28\]\[2\] _05104_ _05105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12324_ _01004_ net526 u_cpu.cpu.ctrl.o_ibus_adr\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06465__I3 u_cpu.rf_ram.memory\[23\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11817__CLK net478 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06870__I0 u_cpu.rf_ram.memory\[104\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12255_ _00938_ net103 u_cpu.rf_ram.memory\[31\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xu_scanchain_local.scan_flop\[35\] u_scanchain_local.module_data_in\[34\] net549 u_arbiter.i_wb_cpu_dbus_dat\[29\]
+ net16 u_scanchain_local.module_data_in\[35\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_29_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11206_ u_cpu.rf_ram.memory\[24\]\[5\] _05493_ _05497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09564__A2 _04312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12186_ _00869_ net497 u_arbiter.i_wb_cpu_dbus_dat\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11137_ _02757_ _05454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_122_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09316__A2 _04143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06202__I _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11068_ u_cpu.rf_ram.memory\[88\]\[0\] _05405_ _05406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10019_ u_cpu.cpu.immdec.imm30_25\[5\] _04672_ _04714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10331__B1 _04931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07878__A2 _03230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout261_I net262 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10882__A1 _05268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout359_I net366 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout526_I net527 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07230_ _02763_ _02792_ _02799_ _00038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11347__CLK net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07161_ _02733_ _02740_ _02742_ _00026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_125_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09252__A1 _04072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06093__B _01709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06112_ _01673_ _01729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_118_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07092_ _02613_ _02616_ _02682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05813__A1 _01456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06861__I0 u_cpu.rf_ram.memory\[36\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06043_ _01659_ _01660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09004__A1 u_cpu.rf_ram.memory\[125\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08799__I _03815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout205 net207 net205 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_114_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07566__A1 _02996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout216 net219 net216 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_134_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09802_ _04431_ _04442_ _04522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06613__I0 u_cpu.rf_ram.memory\[124\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout227 net228 net227 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_86_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout238 net240 net238 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07994_ _03252_ _03312_ _03314_ _00287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout249 net255 net249 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_86_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09307__A2 _04142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09733_ _04416_ _04418_ _04458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06945_ _01408_ _02553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06112__I _01673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07869__A2 _03233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09664_ u_cpu.rf_ram.memory\[113\]\[5\] _04388_ _04392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06876_ _02479_ _02481_ _02483_ _02485_ _01606_ _02486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__10322__B1 _04931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05951__I _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05827_ u_arbiter.i_wb_cpu_dbus_adr\[6\] _01461_ _01470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08615_ _03678_ _03700_ _03707_ _00515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_76_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09595_ _04311_ _04347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12122__CLK net406 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06541__A2 _02146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05758_ _01408_ _01409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08546_ _03600_ _03655_ _03662_ _00491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08039__I _03070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08477_ _03620_ _03622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07097__A3 _02682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09491__A1 _04251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08294__A2 _03488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07428_ _02937_ _02938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_91_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07359_ _02886_ _00080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09794__A2 _04395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10370_ u_cpu.rf_ram.memory\[109\]\[0\] _04962_ _04963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06152__S1 _01768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09029_ _03916_ _03959_ _03967_ _00669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07319__S _02852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12040_ _00723_ net285 u_cpu.rf_ram.memory\[90\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07557__A1 _02987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06604__I0 u_cpu.rf_ram.memory\[108\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06022__I _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07309__A1 _02804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11105__A2 _02572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06957__I _02564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06907__I1 u_cpu.rf_ram.memory\[137\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10864__A1 u_cpu.rf_ram.memory\[108\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11824_ _00520_ net149 u_cpu.rf_ram.memory\[14\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12615__CLK net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11755_ _00451_ net491 u_cpu.rf_ram.memory\[142\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09482__A1 _04242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08285__A2 _03495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07788__I _03180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06906__B _01404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10706_ u_cpu.rf_ram.memory\[104\]\[1\] _05177_ _05179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11686_ _00390_ net299 u_cpu.rf_ram.memory\[57\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06391__S1 _01892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08037__A2 _03338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09234__A1 _04074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10637_ _05130_ _05132_ _05134_ _01111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_70_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10919__A2 _03034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10568_ _05055_ _05085_ _05093_ _01083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07796__A1 _03186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12307_ _00987_ net492 u_cpu.cpu.ctrl.o_ibus_adr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06843__I0 u_cpu.rf_ram.memory\[28\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10499_ _04823_ _05051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_64_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12238_ _00921_ net341 u_cpu.cpu.immdec.imm19_12_20\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12169_ _00852_ net385 u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout476_I net538 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput5 io_in[4] net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_06730_ _02322_ _02341_ _01404_ _02342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_76_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06661_ _01786_ _02272_ _01795_ _02273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10855__A1 _05268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07720__A1 _03119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08400_ _02866_ _03572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_18_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06374__I2 u_cpu.rf_ram.memory\[46\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09380_ _02866_ _04196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_75_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12295__CLK net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06592_ _02198_ _02200_ _02202_ _02204_ _01681_ _02205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_33_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08331_ u_cpu.rf_ram.memory\[54\]\[2\] _03529_ _03530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08276__A2 _03488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11214__S _05501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06287__A1 _01735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10083__A2 _04572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08262_ _03419_ _03474_ _03481_ _00388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07213_ u_cpu.cpu.immdec.imm11_7\[4\] _02787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_140_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09225__A1 u_cpu.rf_ram.memory\[92\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08193_ _03405_ _03439_ _03441_ _00359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07144_ u_cpu.rf_ram_if.genblk1.wtrig0_r _02726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_101_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07075_ u_cpu.rf_ram_if.rdata0\[6\] _02665_ _02669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06026_ u_cpu.rf_ram.memory\[24\]\[0\] u_cpu.rf_ram.memory\[25\]\[0\] u_cpu.rf_ram.memory\[26\]\[0\]
+ u_cpu.rf_ram.memory\[27\]\[0\] _01640_ _01642_ _01643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_126_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07539__A1 _02992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08200__A2 _03439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07977_ u_cpu.rf_ram.memory\[68\]\[2\] _03303_ _03304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09716_ _03113_ u_arbiter.i_wb_cpu_rdt\[15\] _04440_ _04441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_5_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06928_ u_arbiter.i_wb_cpu_dbus_we _02535_ _02536_ _02537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_67_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11512__CLK net319 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09700__A2 _04310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10846__A1 u_cpu.rf_ram.memory\[83\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09647_ _04378_ _04322_ _04329_ _04380_ _04381_ _00874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_71_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06859_ u_cpu.rf_ram.memory\[44\]\[7\] u_cpu.rf_ram.memory\[45\]\[7\] u_cpu.rf_ram.memory\[46\]\[7\]
+ u_cpu.rf_ram.memory\[47\]\[7\] _01721_ _01624_ _02469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07711__A1 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06514__A2 _02121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09578_ u_arbiter.i_wb_cpu_rdt\[8\] _04334_ _04331_ u_arbiter.i_wb_cpu_dbus_dat\[8\]
+ _04335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08529_ u_cpu.rf_ram.memory\[72\]\[6\] _03647_ _03652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11662__CLK net182 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08511__I0 _03576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11540_ _00244_ net249 u_cpu.rf_ram.memory\[77\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10248__B _02691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08019__A2 _03324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11471_ _00175_ net346 u_cpu.rf_ram.memory\[50\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10422_ _04991_ _01039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11023__A1 u_cpu.rf_ram.memory\[86\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12018__CLK net450 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06017__I _01633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10353_ _04949_ _01012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_30_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10284_ _04908_ _04909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12168__CLK net387 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12023_ _00706_ net495 u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09772__B _04494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09063__I _03990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11807_ _00503_ net370 u_cpu.rf_ram.memory\[70\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08258__A2 _03473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10065__A2 _04456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11738_ _00442_ net152 u_cpu.rf_ram.memory\[15\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06364__S1 _01660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09207__A1 _02557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout224_I net228 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11669_ _00373_ net142 u_cpu.rf_ram.memory\[5\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11014__A1 _05354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06992__A2 _01408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07900_ _03227_ _02982_ _03253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08880_ _03560_ u_cpu.rf_ram.memory\[12\]\[0\] _03872_ _03873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_44_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11535__CLK net250 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08194__A1 u_cpu.rf_ram.memory\[19\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06044__I1 u_cpu.rf_ram.memory\[49\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09930__A2 _04629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07831_ _03193_ _03204_ _03211_ _00227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07941__A1 _03264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06595__I2 u_cpu.rf_ram.memory\[46\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07762_ u_cpu.rf_ram.memory\[17\]\[7\] _03153_ _03164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09501_ u_cpu.rf_ram.memory\[33\]\[1\] _04271_ _04273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06713_ u_cpu.rf_ram.memory\[88\]\[5\] u_cpu.rf_ram.memory\[89\]\[5\] u_cpu.rf_ram.memory\[90\]\[5\]
+ u_cpu.rf_ram.memory\[91\]\[5\] _02029_ _01742_ _02325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_53_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07693_ _03114_ _03115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_25_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06644_ _01825_ _02256_ _02257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09432_ _04140_ _04226_ _04228_ _00812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06052__S0 _01639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06898__I3 u_cpu.rf_ram.memory\[71\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09363_ _02845_ _04184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06575_ u_cpu.rf_ram.memory\[20\]\[4\] u_cpu.rf_ram.memory\[21\]\[4\] u_cpu.rf_ram.memory\[22\]\[4\]
+ u_cpu.rf_ram.memory\[23\]\[4\] _01849_ _01965_ _02188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_107_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10056__A2 _02530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08314_ _03498_ _03513_ _03519_ _00402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09997__A2 _04690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09294_ _04074_ _04130_ _04139_ _00763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08245_ u_cpu.rf_ram.memory\[58\]\[7\] _03460_ _03471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11005__A1 _05300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06680__A1 _02285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09749__A2 _04472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08176_ _03426_ _03431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07127_ u_cpu.rf_ram_if.genblk1.wtrig0_r _01387_ _02709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12310__CLK net524 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09148__I _04044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07058_ _02646_ u_cpu.rf_ram_if.rdata1\[5\] _02659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08052__I _03083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06983__A2 _02589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06009_ u_cpu.rf_ram.memory\[16\]\[0\] u_cpu.rf_ram.memory\[17\]\[0\] u_cpu.rf_ram.memory\[18\]\[0\]
+ u_cpu.rf_ram.memory\[19\]\[0\] _01622_ _01625_ _01626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_27_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12460__CLK net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09921__A2 _04398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07932__A1 _03252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06586__I2 u_cpu.rf_ram.memory\[50\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10819__A1 _05206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09685__A1 _01440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08488__A2 _03621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10971_ u_cpu.rf_ram.memory\[85\]\[5\] _05340_ _05344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10295__A2 _04915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07160__A2 _02741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12641_ _01320_ net64 u_cpu.rf_ram.memory\[24\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09437__A1 _04147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10047__A2 _04636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[60\]_SE net554 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12572_ _01251_ net200 u_cpu.rf_ram.memory\[86\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07999__A1 _03259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11408__CLK net224 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11523_ _00227_ net431 u_cpu.rf_ram.memory\[129\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08660__A2 _02940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06970__I _01387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11454_ _00158_ net334 u_cpu.rf_ram.memory\[48\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10405_ _02723_ _02850_ _04982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__10492__I _04816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11385_ _00089_ net217 u_cpu.rf_ram.memory\[80\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11558__CLK net250 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09058__I _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06423__A1 _02028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06274__I1 u_cpu.rf_ram.memory\[109\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10336_ u_cpu.cpu.ctrl.o_ibus_adr\[21\] _04936_ _04938_ u_cpu.cpu.ctrl.o_ibus_adr\[22\]
+ _04940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_106_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06974__A2 _02547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10267_ _04893_ _04898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08897__I _03881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12006_ _00689_ net409 u_cpu.rf_ram.memory\[37\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09912__A2 _04548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10198_ u_arbiter.i_wb_cpu_dbus_adr\[9\] u_arbiter.i_wb_cpu_dbus_adr\[8\] _04855_
+ _04857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07923__A1 _03268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06577__I2 u_cpu.rf_ram.memory\[18\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06282__S0 _01729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06210__I _01788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout174_I net176 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08479__A2 _03621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10286__A2 _04907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout341_I net344 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10667__I _05150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09428__A1 _02937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout439_I net440 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11235__A1 u_cpu.rf_ram.memory\[98\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06360_ _01857_ _01974_ _01859_ _01975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09979__A2 _04566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08100__A1 _03380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06291_ _01904_ _01906_ _01744_ _01907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07976__I _03298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08030_ _03059_ _03335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09600__A1 u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12483__CLK net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09981_ _04420_ _04492_ _04676_ _04678_ _04679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__06965__A2 _02572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08932_ _02756_ _03906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout87_I net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08167__A1 _03423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09903__A2 _04432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08863_ _03819_ _03859_ _03862_ _00608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07914__A1 _03262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07814_ u_cpu.rf_ram.memory\[119\]\[7\] _03182_ _03200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08794_ _03813_ _03816_ _03818_ _00583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07216__I _02789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07390__A2 _02901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06120__I _01687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07745_ _03153_ _03154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09667__A1 _04253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10277__A2 _04895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07676_ _03104_ _00179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09415_ u_cpu.rf_ram.memory\[112\]\[2\] _04217_ _04218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09419__A1 u_cpu.rf_ram.memory\[112\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06627_ u_cpu.rf_ram.memory\[80\]\[4\] u_cpu.rf_ram.memory\[81\]\[4\] u_cpu.rf_ram.memory\[82\]\[4\]
+ u_cpu.rf_ram.memory\[83\]\[4\] _01651_ _02033_ _02240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_90_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10029__A2 _04549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09346_ u_cpu.rf_ram.memory\[121\]\[0\] _04174_ _04175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06558_ u_cpu.rf_ram.memory\[128\]\[3\] u_cpu.rf_ram.memory\[129\]\[3\] u_cpu.rf_ram.memory\[130\]\[3\]
+ u_cpu.rf_ram.memory\[131\]\[3\] _01826_ _01827_ _02172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_90_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09277_ _04128_ _04130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06489_ _01687_ _02103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_103_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08228_ _03460_ _03461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11700__CLK net425 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08159_ _03080_ _03419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09807__S _04417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11170_ u_cpu.rf_ram.memory\[26\]\[7\] _05464_ _05475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10121_ u_cpu.cpu.genblk3.csr.timer_irq_r _04804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_79_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11850__CLK net508 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08158__A1 _03417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07327__S _02852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10052_ u_cpu.cpu.immdec.imm19_12_20\[2\] _04743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_7_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[8\]_SI u_arbiter.i_wb_cpu_dbus_dat\[2\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06264__S0 _01692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12206__CLK net383 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06030__I _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10268__A2 _04898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10954_ _05333_ _01229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07133__A2 _02714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10885_ _05288_ _05293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_43_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06892__A1 _02147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12624_ _01303_ net57 u_cpu.rf_ram.memory\[26\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06319__S1 _01799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[65\] u_scanchain_local.module_data_in\[64\] net554 u_arbiter.o_wb_cpu_adr\[27\]
+ net22 u_scanchain_local.module_data_in\[65\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_12_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12555_ _01234_ net211 u_cpu.rf_ram.memory\[85\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09830__A1 _04427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06914__B _01644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11380__CLK net176 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11506_ _00210_ net326 u_cpu.rf_ram.memory\[40\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12486_ _01165_ net39 u_cpu.rf_ram.memory\[105\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11437_ _00141_ net324 u_cpu.rf_ram.memory\[41\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11368_ _00072_ net134 u_cpu.rf_ram.memory\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09944__C _04526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06947__A2 _02549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10319_ _01502_ _04929_ _04924_ u_cpu.cpu.ctrl.o_ibus_adr\[15\] _04930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11299_ _02899_ _05547_ _05552_ _01355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout291_I net294 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout389_I net391 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09897__A1 _04403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05860_ u_arbiter.i_wb_cpu_dbus_adr\[12\] _01481_ _01497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09960__B _04427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10598__S _05111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05791_ _01437_ _01438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_81_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout556_I net557 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10259__A2 _04888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07530_ _03006_ _03008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_78_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06558__S1 _01827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07461_ u_cpu.rf_ram.memory\[46\]\[3\] _02958_ _02960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06183__I0 u_cpu.rf_ram.memory\[72\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08872__A2 _03860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09200_ _02549_ _04079_ _04080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06722__I2 u_cpu.rf_ram.memory\[70\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06412_ u_cpu.rf_ram.memory\[92\]\[2\] u_cpu.rf_ram.memory\[93\]\[2\] u_cpu.rf_ram.memory\[94\]\[2\]
+ u_cpu.rf_ram.memory\[95\]\[2\] _01762_ _01915_ _02027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_72_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07392_ _02772_ _02912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09131_ _04031_ _04030_ _04033_ _00705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06343_ _01398_ _01958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_17_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11222__S _05501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09062_ _03990_ _03991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06274_ u_cpu.rf_ram.memory\[108\]\[1\] u_cpu.rf_ram.memory\[109\]\[1\] u_cpu.rf_ram.memory\[110\]\[1\]
+ u_cpu.rf_ram.memory\[111\]\[1\] _01716_ _01717_ _01890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_50_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07683__I0 _02867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08013_ u_cpu.rf_ram.memory\[66\]\[0\] _03325_ _03326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09585__B1 _04331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09964_ _04585_ _04663_ _04664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_131_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08915_ _03832_ _03883_ _03892_ _00630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09895_ u_arbiter.i_wb_cpu_rdt\[5\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[5\]
+ _01440_ _04601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09888__A1 _04251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08846_ _03821_ _03847_ _03852_ _00601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08560__A1 u_cpu.rf_ram.memory\[71\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08777_ _03752_ _03802_ _03807_ _00577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_2_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12379__CLK net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05989_ _01605_ _01606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_2827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07728_ _03060_ _03142_ _03144_ _00191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08312__A1 _03494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07659_ u_cpu.rf_ram.memory\[50\]\[2\] _03094_ _03095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08863__A2 _03859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10670_ u_cpu.rf_ram.memory\[102\]\[3\] _05155_ _05157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09329_ _04145_ _04161_ _04164_ _00773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09812__A1 _02557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08615__A2 _03700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06734__B _01628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06626__A1 _01740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12340_ _01020_ net165 u_cpu.rf_ram.memory\[109\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12271_ _00954_ net530 u_arbiter.i_wb_cpu_dbus_adr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11222_ _02863_ u_cpu.rf_ram.memory\[0\]\[4\] _05501_ _05506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06025__I _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09040__A2 _03973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10770__I _05219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11153_ _05464_ _05465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_66_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10104_ u_cpu.cpu.immdec.imm19_12_20\[7\] _04739_ _04790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11084_ _05365_ _05405_ _05414_ _01278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09879__A1 _04242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10035_ _04416_ _04724_ _04728_ _04729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_103_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08551__A1 u_cpu.rf_ram.memory\[73\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06401__I1 u_cpu.rf_ram.memory\[125\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10211__S _04861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11986_ _00676_ net439 u_cpu.rf_ram.memory\[123\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08303__A1 _02877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10110__A1 _04397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10937_ u_cpu.rf_ram.memory\[59\]\[7\] _05313_ _05324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08854__A2 _03848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06865__B2 _02474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10868_ _05280_ _05270_ _05281_ _01195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12607_ _01286_ net380 u_cpu.cpu.genblk3.csr.mstatus_mie vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11896__CLK net459 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout137_I net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08606__A2 _03700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10799_ u_cpu.rf_ram.memory\[106\]\[3\] _05236_ _05238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12538_ _01217_ net279 u_cpu.rf_ram.memory\[59\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06468__I1 u_cpu.rf_ram.memory\[17\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06093__A2 _01708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout304_I net305 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07290__A1 u_cpu.rf_ram.memory\[20\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12469_ _01148_ net46 u_cpu.rf_ram.memory\[99\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09031__A2 _03959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10680__I _04958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06476__S0 _01863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout409 net412 net409 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_119_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08790__A1 _02786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07593__A2 _03005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06961_ u_cpu.cpu.bufreg2.i_cnt_done _02569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08700_ u_cpu.rf_ram.memory\[137\]\[5\] _03753_ _03760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05912_ u_cpu.cpu.ctrl.o_ibus_adr\[24\] _01537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_95_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06228__S0 _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09680_ _01439_ _04405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06892_ _02147_ _02501_ _02502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08542__A1 _03595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08631_ _03716_ _00522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05843_ _01473_ _01480_ _01482_ u_arbiter.o_wb_cpu_adr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08562_ _03493_ _03673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05774_ u_cpu.cpu.immdec.imm24_20\[2\] _01389_ _01425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09098__A2 _04004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12671__CLK net288 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07513_ u_cpu.rf_ram.memory\[44\]\[4\] _02990_ _02995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08493_ u_cpu.rf_ram.memory\[140\]\[7\] _03620_ _03631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08845__A2 _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09893__I1 u_arbiter.i_wb_cpu_rdt\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout16 net18 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout27 net32 net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06856__A1 _02459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10652__A2 _05138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout38 net42 net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_50_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07444_ _02907_ _02942_ _02949_ _00102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout49 net50 net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_11_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07375_ _02751_ _02899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05949__I _01565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09114_ _03982_ _04015_ _04022_ _00699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06326_ _01815_ _01942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06703__S1 _01905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09045_ _03977_ _03972_ _03979_ _00673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06257_ _01678_ _01873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06084__A2 _01700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06188_ _01418_ _01805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09022__A2 _03962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07584__A2 _03036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08781__A1 _03757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09947_ u_cpu.cpu.immdec.imm24_20\[3\] _04629_ _04649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09878_ u_cpu.rf_ram.memory\[114\]\[1\] _04589_ _04591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11769__CLK net481 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08533__A1 _03272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08829_ u_cpu.rf_ram.memory\[132\]\[4\] _03839_ _03842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10340__B2 _01537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11840_ _00536_ net421 u_cpu.rf_ram.memory\[39\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10891__A2 _05289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09089__A2 _04007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11771_ _00467_ net491 u_cpu.rf_ram.memory\[140\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06147__I0 u_cpu.rf_ram.memory\[92\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08836__A2 _03836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10722_ _05187_ _05188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10643__A2 _05138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10653_ _05144_ _05133_ _05145_ _01116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10584_ _05099_ _05104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12323_ _01003_ net526 u_cpu.cpu.ctrl.o_ibus_adr\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07272__A1 _02763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05822__A2 _01461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12254_ _00937_ net97 u_cpu.rf_ram.memory\[31\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10159__A1 u_cpu.rf_ram.memory\[32\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11205_ _05456_ _05489_ _05496_ _01317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06458__S0 _01959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_scanchain_local.scan_flop\[28\] u_arbiter.i_wb_cpu_rdt\[25\] net547 u_arbiter.i_wb_cpu_dbus_dat\[22\]
+ net17 u_arbiter.i_wb_cpu_rdt\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
X_12185_ _00868_ net390 u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08772__A1 _03745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11136_ _05451_ _05446_ _05453_ _01291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10005__I _04505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11067_ _05403_ _05405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_42_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08524__A1 _03598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12694__CLK net379 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10018_ _04499_ _04706_ _04712_ _04395_ _04713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_77_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05889__A2 _01516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10882__A2 _05289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07314__I _02854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout254_I net255 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08827__A2 _03839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11969_ _00665_ net446 u_cpu.rf_ram.memory\[124\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout421_I net423 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout519_I net520 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07160_ u_cpu.rf_ram.memory\[82\]\[0\] _02741_ _02742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09252__A2 _04106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06111_ _01595_ _01728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07263__A1 _02740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07091_ _02676_ _02680_ _02681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06042_ _01658_ _01659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09004__A2 _03950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07015__A1 _02553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10945__I0 _04190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout206 net207 net206 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_119_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09801_ _04514_ _04423_ _04506_ _04521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout217 net219 net217 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__08763__A1 _03759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06613__I1 u_cpu.rf_ram.memory\[125\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout228 net229 net228 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__11911__CLK net457 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07993_ u_cpu.rf_ram.memory\[67\]\[0\] _03313_ _03314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout239 net240 net239 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__10570__A1 _05057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09732_ _04456_ _04457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06944_ _02530_ _02533_ _02552_ _00021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09663_ _04249_ _04384_ _04391_ _00880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06875_ _01720_ _02484_ _01663_ _02485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_39_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08614_ u_cpu.rf_ram.memory\[143\]\[4\] _03704_ _03707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05826_ _01434_ _01468_ _01469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09594_ u_arbiter.i_wb_cpu_dbus_dat\[14\] _04338_ _04346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10873__A2 _05276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07224__I _02791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08545_ u_cpu.rf_ram.memory\[73\]\[4\] _03659_ _03662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05757_ u_cpu.cpu.csr_d_sel _01408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06829__A1 _01406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12417__CLK net357 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08476_ _03620_ _03621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07427_ _02721_ _02936_ _02937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_50_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08055__I _03086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07358_ _02870_ u_cpu.rf_ram.memory\[7\]\[6\] _02878_ _02886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_13_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09243__A2 _04109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06309_ _01426_ _01925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07254__A1 _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11441__CLK net325 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11050__A2 _05393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12567__CLK net163 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07289_ _02832_ _02837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09028_ u_cpu.rf_ram.memory\[124\]\[6\] _03962_ _03967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[17\]_SE net542 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08754__A1 _03750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10561__A1 u_cpu.rf_ram.memory\[96\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07309__A2 _02850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07335__S _02851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06368__I0 u_cpu.rf_ram.memory\[56\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06907__I2 u_cpu.rf_ram.memory\[138\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10864__A2 _05276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11823_ _00519_ net136 u_cpu.rf_ram.memory\[14\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08809__A2 _03822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12097__CLK net410 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11754_ _00450_ net490 u_cpu.rf_ram.memory\[142\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09482__A2 _04258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10705_ _05130_ _05176_ _05178_ _01135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07493__A1 _02916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11685_ _00389_ net287 u_cpu.rf_ram.memory\[57\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06194__B _01810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10636_ u_cpu.rf_ram.memory\[101\]\[0\] _05133_ _05134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_u_scanchain_local.scan_flop\[31\]_D u_arbiter.i_wb_cpu_rdt\[28\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07245__A1 _02746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11041__A2 _05384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10567_ u_cpu.rf_ram.memory\[96\]\[6\] _05088_ _05093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12306_ _00986_ net503 u_cpu.cpu.ctrl.o_ibus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06843__I1 u_cpu.rf_ram.memory\[29\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11934__CLK net333 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10498_ _05049_ _05041_ _05050_ _01056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_12237_ _00920_ net359 u_cpu.cpu.csr_imm vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08745__A1 _03761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06213__I _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12168_ _00851_ net387 u_arbiter.i_wb_cpu_dbus_dat\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11119_ _05438_ _05439_ _05440_ _05441_ _01286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__06220__A2 _01836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12099_ _00782_ net448 u_cpu.rf_ram.memory\[121\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout371_I net372 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout469_I net472 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06660_ u_cpu.rf_ram.memory\[0\]\[5\] u_cpu.rf_ram.memory\[1\]\[5\] u_cpu.rf_ram.memory\[2\]\[5\]
+ u_cpu.rf_ram.memory\[3\]\[5\] _02074_ _01585_ _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10855__A2 _05270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06591_ _02098_ _02203_ _01873_ _02204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08330_ _03524_ _03529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_75_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06816__C _02050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06287__A2 _01902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08261_ u_cpu.rf_ram.memory\[57\]\[5\] _03477_ _03481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11464__CLK net226 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06531__I0 u_cpu.rf_ram.memory\[88\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07212_ _02785_ _02786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_14_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[22\]_D u_arbiter.i_wb_cpu_rdt\[19\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08192_ u_cpu.rf_ram.memory\[19\]\[0\] _03440_ _03441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09225__A2 _04097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07236__A1 _02778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07143_ u_cpu.cpu.immdec.imm11_7\[2\] _02724_ _02725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07074_ _02662_ _02656_ _02668_ _00012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05798__A1 _01443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06025_ _01641_ _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08736__A1 u_cpu.rf_ram.memory\[136\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07219__I _02791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07539__A2 _03007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06123__I _01671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10543__A1 u_cpu.rf_ram.memory\[95\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07976_ _03298_ _03303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_75_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09715_ _01438_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\] _04440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_142_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06927_ u_cpu.cpu.decode.opcode\[2\] u_cpu.cpu.decode.opcode\[1\] u_cpu.cpu.decode.opcode\[0\]
+ _02536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_68_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09161__A1 u_cpu.rf_ram.memory\[91\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09646_ u_arbiter.i_wb_cpu_rdt\[30\] _04300_ _04381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10846__A2 _05261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06858_ _01772_ _02467_ _02468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07711__A2 _01450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05809_ _01451_ _01455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09577_ _04311_ _04334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11807__CLK net370 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06789_ u_cpu.rf_ram.memory\[124\]\[6\] u_cpu.rf_ram.memory\[125\]\[6\] u_cpu.rf_ram.memory\[126\]\[6\]
+ u_cpu.rf_ram.memory\[127\]\[6\] _02015_ _01774_ _02400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_93_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08528_ _03602_ _03644_ _03651_ _00484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_19_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06278__A2 _01893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08459_ _03588_ _03609_ _03611_ _00455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[13\]_D u_arbiter.i_wb_cpu_rdt\[10\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_11470_ _00174_ net347 u_cpu.rf_ram.memory\[50\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11957__CLK net441 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10421_ _04200_ u_cpu.rf_ram.memory\[2\]\[7\] _04982_ _04991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07227__A1 u_cpu.rf_ram.memory\[21\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07778__A2 _03172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10352_ u_cpu.cpu.ctrl.o_ibus_adr\[28\] _04943_ _04945_ u_cpu.cpu.ctrl.o_ibus_adr\[29\]
+ _04949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_3_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10782__A1 _05211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06450__A2 _02064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10283_ net2 _02696_ _04908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08727__A1 _03763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12022_ _00705_ net482 u_cpu.cpu.mem_bytecnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06033__I _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11337__CLK net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09152__A1 u_cpu.rf_ram.memory\[91\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11487__CLK net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06917__B _02526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11806_ _00502_ net347 u_cpu.rf_ram.memory\[71\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09455__A2 _04240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07466__A1 _02910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11737_ _00441_ net149 u_cpu.rf_ram.memory\[15\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11262__A2 _05527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06208__I _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08624__S _03712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11668_ _00372_ net122 u_cpu.rf_ram.memory\[5\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10619_ _03116_ _05123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__11014__A2 _05368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout217_I net219 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11599_ _00303_ net244 u_cpu.rf_ram.memory\[65\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10773__A1 _05199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12112__CLK net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08718__A1 u_cpu.rf_ram.memory\[49\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09915__B1 _04523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10525__A1 u_cpu.rf_ram.memory\[94\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08194__A2 _03440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07830_ u_cpu.rf_ram.memory\[129\]\[4\] _03208_ _03211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06044__I2 u_cpu.rf_ram.memory\[50\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05782__I u_arbiter.i_wb_cpu_ibus_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12262__CLK net491 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[40\]_CLK net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07941__A2 _03274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06595__I3 u_cpu.rf_ram.memory\[47\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07761_ _03084_ _03155_ _03163_ _00205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09500_ _04237_ _04270_ _04272_ _00836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06712_ _01735_ _02323_ _02324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10828__A2 _05244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07692_ _03113_ _03114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_64_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09431_ u_cpu.rf_ram.memory\[122\]\[0\] _04227_ _04228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06643_ u_cpu.rf_ram.memory\[136\]\[4\] u_cpu.rf_ram.memory\[137\]\[4\] u_cpu.rf_ram.memory\[138\]\[4\]
+ u_cpu.rf_ram.memory\[139\]\[4\] _01814_ _01942_ _02256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_24_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout32_I net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09362_ _04158_ _04174_ _04183_ _00787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06574_ _02180_ _02182_ _02184_ _02186_ _01607_ _02187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_21_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09446__A2 _04225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07502__I _02896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08313_ u_cpu.rf_ram.memory\[55\]\[3\] _03517_ _03519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07457__A1 _02897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10056__A3 _04482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11253__A2 _05524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06504__I0 u_cpu.rf_ram.memory\[108\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09293_ u_cpu.rf_ram.memory\[117\]\[7\] _04128_ _04139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08244_ _03421_ _03462_ _03470_ _00381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06118__I _01648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07209__A1 _02708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11005__A2 _03286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08175_ _03410_ _03427_ _03430_ _00352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06680__A2 _02287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05957__I _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06562__B _01419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09429__I _04225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07126_ _01387_ _01395_ u_cpu.rf_ram_if.genblk1.wtrig0_r _02708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10764__A1 u_cpu.rf_ram.memory\[79\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07057_ _02542_ u_cpu.rf_ram.rdata\[5\] _02658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06008_ _01624_ _01625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12605__CLK net378 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10516__A1 u_cpu.rf_ram.memory\[94\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08185__A2 _03431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07932__A2 _03274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07959_ _02861_ u_cpu.rf_ram.memory\[6\]\[3\] _03289_ _03293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_46_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09134__A1 _04034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10970_ _05280_ _05336_ _05343_ _01235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10819__A2 _05245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07145__B1 u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09685__A2 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09629_ _04368_ _04369_ _00868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06499__A2 _02112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12640_ _01319_ net67 u_cpu.rf_ram.memory\[24\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09437__A2 _04226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07448__A1 _02913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12571_ _01250_ net200 u_cpu.rf_ram.memory\[86\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11244__A2 _05515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10452__B1 _04652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07999__A2 _03312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11522_ _00226_ net430 u_cpu.rf_ram.memory\[129\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12135__CLK net436 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11453_ _00157_ net334 u_cpu.rf_ram.memory\[48\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10404_ _04981_ _01031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11384_ _00088_ net217 u_cpu.rf_ram.memory\[80\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06191__C _01807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10335_ _04939_ _01004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06423__A2 _02032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07620__A1 u_cpu.rf_ram.memory\[47\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12285__CLK net505 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10266_ _04814_ _04894_ _04897_ _00977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10507__A1 _05055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[10\] u_arbiter.i_wb_cpu_rdt\[7\] net544 u_arbiter.i_wb_cpu_dbus_dat\[4\]
+ net12 u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
X_12005_ _00688_ net408 u_cpu.rf_ram.memory\[37\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06026__I2 u_cpu.rf_ram.memory\[26\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10197_ _04856_ _00949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07923__A2 _03255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06577__I3 u_cpu.rf_ram.memory\[19\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06282__S1 _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout167_I net172 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07322__I _02860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09428__A2 _04224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11235__A2 _05512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09979__A3 _04659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout334_I net335 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08100__A2 _03062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06290_ u_cpu.rf_ram.memory\[120\]\[1\] u_cpu.rf_ram.memory\[121\]\[1\] u_cpu.rf_ram.memory\[122\]\[1\]
+ u_cpu.rf_ram.memory\[123\]\[1\] _01741_ _01905_ _01906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_15_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout501_I net502 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10683__I _05163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05777__I _01427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08939__A1 _03910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08153__I _03074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11502__CLK net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12628__CLK net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10746__A1 _05199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09600__A2 _04338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09980_ _04545_ _04677_ _04678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07992__I _03311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08931_ _03903_ _03896_ _03905_ _00633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11652__CLK net220 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08167__A2 _03408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08411__I0 _03560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08862_ u_cpu.rf_ram.memory\[130\]\[1\] _03860_ _03862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11171__A1 _05462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07914__A2 _03254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07813_ _03086_ _03199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_29_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08793_ u_cpu.rf_ram.memory\[133\]\[0\] _03817_ _03818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09116__A1 _03984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07744_ _02790_ _02804_ _03153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09667__A2 _04385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07675_ _02855_ u_cpu.rf_ram.memory\[4\]\[1\] _03102_ _03104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_52_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06557__B _01823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09414_ _04212_ _04217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06626_ _01740_ _02238_ _02031_ _02239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_41_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09345_ _04172_ _04174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10029__A3 _04434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06557_ _01819_ _02170_ _01823_ _02171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09276_ _04128_ _04129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06102__A1 _01715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06488_ _02091_ _02094_ _02097_ _02101_ _01681_ _02102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__10985__A1 _05352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08227_ _02937_ _03425_ _03460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08158_ _03417_ _03407_ _03418_ _00347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07109_ _01431_ u_cpu.cpu.ctrl.pc_plus_4_cy_r _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07602__A1 _02989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08089_ u_cpu.rf_ram.memory\[29\]\[3\] _03373_ _03375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10120_ _04467_ _04619_ _04801_ _04803_ _00925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__06956__A3 u_cpu.cpu.mem_bytecnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08158__A2 _03407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10051_ _04741_ _04738_ _04742_ _04531_ _00917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_88_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05916__A1 _01524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06264__S1 _01879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09107__A1 _03975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09658__A2 _04388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07669__A1 u_cpu.rf_ram.memory\[50\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10953_ _04198_ u_cpu.rf_ram.memory\[10\]\[6\] _05325_ _05333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_16_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10884_ _05273_ _05289_ _05292_ _01200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12623_ _01302_ net52 u_cpu.rf_ram.memory\[26\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06892__A2 _02501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12554_ _01233_ net212 u_cpu.rf_ram.memory\[85\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08094__A1 _03349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11525__CLK net430 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10976__A1 _05286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09830__A2 _04546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11505_ _00209_ net302 u_cpu.rf_ram.memory\[40\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06644__A2 _02256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[58\] u_scanchain_local.module_data_in\[57\] net562 u_arbiter.o_wb_cpu_adr\[20\]
+ net30 u_scanchain_local.module_data_in\[58\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__10209__S _04861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12485_ _01164_ net41 u_cpu.rf_ram.memory\[105\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11436_ _00140_ net327 u_cpu.rf_ram.memory\[41\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11675__CLK net325 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11367_ _00071_ net123 u_cpu.rf_ram.memory\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10318_ _04905_ _04929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11298_ u_cpu.rf_ram.memory\[23\]\[2\] _05551_ _05552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10249_ _02675_ _02627_ _02686_ _02688_ _04885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_67_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09897__A2 _04602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10200__I0 u_arbiter.i_wb_cpu_dbus_adr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout284_I net285 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05790_ u_cpu.cpu.genblk1.align.ctrl_misal _01437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_94_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09649__A2 _04322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06580__A1 _01630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout451_I net452 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout549_I net550 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12300__CLK net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07460_ _02900_ _02954_ _02959_ _00108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06183__I1 u_cpu.rf_ram.memory\[73\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06411_ _01565_ _02026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06722__I3 u_cpu.rf_ram.memory\[71\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11208__A2 _05493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07391_ _02910_ _02894_ _02911_ _00087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09130_ _04031_ _04030_ _04032_ _04033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06342_ _01580_ _01956_ _01588_ _01957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08085__A1 _03340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09061_ _03018_ _03286_ _03990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06635__A2 _02247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07832__A1 u_cpu.rf_ram.memory\[129\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06273_ _01566_ _01848_ _01861_ _01888_ _01889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__08880__I0 _03560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08012_ _03323_ _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10719__A1 u_cpu.rf_ram.memory\[104\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09585__A1 u_arbiter.i_wb_cpu_rdt\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08632__I0 _03570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09963_ _04528_ _04484_ _04486_ _04658_ _04662_ _04663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_98_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09337__A1 u_cpu.rf_ram.memory\[118\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08914_ u_cpu.rf_ram.memory\[22\]\[7\] _03881_ _03892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09894_ _04499_ _04599_ _04600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11144__A1 u_cpu.rf_ram.memory\[27\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[50\]_SE net558 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10081__C _04768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06131__I _01652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08845_ u_cpu.rf_ram.memory\[131\]\[2\] _03851_ _03852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08776_ u_cpu.rf_ram.memory\[134\]\[2\] _03806_ _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05988_ _01424_ _01425_ _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06571__A1 _01958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05970__I _01417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07727_ u_cpu.rf_ram.memory\[16\]\[0\] _03143_ _03144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08312__A2 _03513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11548__CLK net339 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07658_ _03089_ _03094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06323__A1 _01928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06609_ _02008_ _02221_ _02222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06713__I3 u_cpu.rf_ram.memory\[91\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07589_ u_cpu.rf_ram.memory\[43\]\[6\] _03040_ _03045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09328_ u_cpu.rf_ram.memory\[118\]\[1\] _04162_ _04164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08076__A1 u_cpu.rf_ram.memory\[64\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09812__A2 _04396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11698__CLK net452 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09259_ _04056_ _04117_ _04119_ _00748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07823__A1 u_cpu.rf_ram.memory\[129\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12270_ _00953_ net530 u_arbiter.i_wb_cpu_dbus_adr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06306__I _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11221_ _05505_ _01324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08379__A2 _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11152_ _05098_ _02938_ _05464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09328__A1 u_cpu.rf_ram.memory\[118\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10103_ u_cpu.cpu.immdec.imm19_12_20\[8\] _04395_ _04789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11083_ u_cpu.rf_ram.memory\[88\]\[7\] _05403_ _05414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10034_ _04721_ _04710_ _04725_ _04727_ _04474_ _04728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__06041__I u_cpu.raddr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06237__S1 _01625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[3\] u_arbiter.i_wb_cpu_rdt\[0\] net547 u_arbiter.i_wb_cpu_dbus_sel\[1\]
+ net17 u_arbiter.i_wb_cpu_rdt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_62_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06562__A1 _02060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11985_ _00675_ net438 u_cpu.rf_ram.memory\[123\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09500__A1 _04237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08303__A2 _03425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10936_ _05284_ _05315_ _05323_ _01221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_90_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12473__CLK net241 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10867_ u_cpu.rf_ram.memory\[108\]\[4\] _05276_ _05281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08067__A1 _03342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12606_ _01285_ net480 u_cpu.cpu.genblk3.csr.mie_mtie vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10798_ _05206_ _05232_ _05237_ _01169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07600__I _03047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12537_ _01216_ net278 u_cpu.rf_ram.memory\[59\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07814__A1 u_cpu.rf_ram.memory\[119\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06468__I2 u_cpu.rf_ram.memory\[18\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08632__S _03712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12468_ _01147_ net46 u_cpu.rf_ram.memory\[99\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07290__A2 _02837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11419_ _00123_ net291 u_cpu.rf_ram.memory\[44\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12399_ _01078_ net44 u_cpu.rf_ram.memory\[96\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10177__A2 _04840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06476__S1 _01653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout499_I net506 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09319__A1 _04156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08790__A2 _03814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09971__B _04667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06960_ u_cpu.cpu.genblk3.csr.mcause3_0\[0\] _02568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input4_I io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05911_ _01453_ _01533_ _01535_ _01536_ u_arbiter.o_wb_cpu_adr\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__06228__S1 _01592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06891_ u_cpu.rf_ram.memory\[80\]\[7\] u_cpu.rf_ram.memory\[81\]\[7\] u_cpu.rf_ram.memory\[82\]\[7\]
+ u_cpu.rf_ram.memory\[83\]\[7\] _01651_ _01653_ _02501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_132_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08630_ _03568_ u_cpu.rf_ram.memory\[14\]\[3\] _03712_ _03716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08542__A2 _03655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05842_ u_arbiter.i_wb_cpu_dbus_adr\[9\] _01481_ _01482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05790__I u_cpu.cpu.genblk1.align.ctrl_misal vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08561_ _03671_ _03668_ _03672_ _00496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05773_ u_cpu.cpu.immdec.imm19_12_20\[6\] _01367_ _01424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07512_ _02906_ _02994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08492_ _03604_ _03622_ _03630_ _00469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06305__A1 _01772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10101__A2 _04786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout17 net18 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07443_ u_cpu.rf_ram.memory\[42\]\[4\] _02946_ _02949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout28 net32 net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__06856__A2 _02461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout39 net42 net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__11840__CLK net421 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08058__A1 _02891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07374_ _02897_ _02893_ _02898_ _00083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout9_I net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09113_ u_cpu.rf_ram.memory\[36\]\[4\] _04019_ _04022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06325_ _01914_ _01940_ _01810_ _01941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07805__A1 u_cpu.rf_ram.memory\[119\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11032__I _05379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06164__S0 _01779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09044_ u_cpu.rf_ram.memory\[123\]\[2\] _03978_ _03979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06256_ u_cpu.rf_ram.memory\[56\]\[1\] u_cpu.rf_ram.memory\[57\]\[1\] u_cpu.rf_ram.memory\[58\]\[1\]
+ u_cpu.rf_ram.memory\[59\]\[1\] _01871_ _01676_ _01872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__11990__CLK net263 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06187_ u_cpu.rf_ram.memory\[76\]\[0\] u_cpu.rf_ram.memory\[77\]\[0\] u_cpu.rf_ram.memory\[78\]\[0\]
+ u_cpu.rf_ram.memory\[79\]\[0\] _01582_ _01803_ _01804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_132_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05965__I _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08781__A2 _03802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09946_ u_cpu.cpu.immdec.imm24_20\[4\] _04572_ _04648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11117__A1 _04952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06792__A1 _01672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09877_ _04237_ _04588_ _04590_ _00895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09730__A1 _04403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08533__A2 _03020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08828_ _03824_ _03835_ _03841_ _00594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11370__CLK net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10340__A2 _04936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08759_ _03755_ _03790_ _03796_ _00570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11770_ _00466_ net490 u_cpu.rf_ram.memory\[140\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08297__A1 u_cpu.rf_ram.memory\[56\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10721_ _03002_ _05162_ _05187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10652_ u_cpu.rf_ram.memory\[101\]\[5\] _05138_ _05145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09797__A1 _04415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10583_ _05044_ _05100_ _05103_ _01088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_12322_ _01002_ net532 u_cpu.cpu.ctrl.o_ibus_adr\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06036__I _01652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07272__A2 _02818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12253_ _00936_ net93 u_cpu.rf_ram.memory\[31\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10159__A2 _04809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11204_ u_cpu.rf_ram.memory\[24\]\[4\] _05493_ _05496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11098__B _02693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12184_ _00867_ net389 u_arbiter.i_wb_cpu_dbus_dat\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06458__S1 _02071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06083__I0 u_cpu.rf_ram.memory\[36\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11135_ u_cpu.rf_ram.memory\[27\]\[2\] _05452_ _05453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08772__A2 _03802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11713__CLK net450 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11066_ _05403_ _05404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_48_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10017_ _04708_ _04711_ _04619_ _04712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08524__A2 _03643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10222__S _04867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05824__B u_cpu.cpu.ctrl.o_ibus_adr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06535__A1 _02147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10331__A2 _04936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05969__S0 _01583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11863__CLK net516 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07335__I0 _02870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11968_ _00664_ net463 u_cpu.rf_ram.memory\[124\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10919_ _03004_ _03034_ _05313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout247_I net248 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11899_ _00595_ net471 u_cpu.rf_ram.memory\[132\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06394__S0 _01621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12219__CLK net318 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07330__I _02866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06110_ _01725_ _01726_ _01727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07090_ u_cpu.cpu.decode.opcode\[1\] _02680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07263__A2 _02818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06041_ u_cpu.raddr\[1\] _01658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_12_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05785__I _01433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07015__A2 _02620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09800_ _04519_ _04520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09960__A1 _04492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08763__A2 _03791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout207 net208 net207 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_113_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout218 net219 net218 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07992_ _03311_ _03313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout229 net230 net229 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_119_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11393__CLK net249 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06774__A1 _01715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09731_ _04450_ _04453_ _04455_ _04456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_06943_ _02530_ _02551_ _02552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11228__S _05500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09662_ u_cpu.rf_ram.memory\[113\]\[4\] _04388_ _04391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06874_ u_cpu.rf_ram.memory\[96\]\[7\] u_cpu.rf_ram.memory\[97\]\[7\] u_cpu.rf_ram.memory\[98\]\[7\]
+ u_cpu.rf_ram.memory\[99\]\[7\] _02125_ _01693_ _02484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA_fanout62_I net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10322__A2 _04929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06526__B2 _02138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07505__I _02899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08613_ _03676_ _03700_ _03706_ _00514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05825_ u_cpu.cpu.ctrl.o_ibus_adr\[6\] _01463_ _01464_ _01468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09593_ _04343_ _04345_ _00856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11027__I _05379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08544_ _03598_ _03655_ _03661_ _00490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05756_ u_cpu.cpu.immdec.imm19_12_20\[5\] u_cpu.rf_ram_if.rtrig0 _01407_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10086__A1 _04738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08475_ _02981_ _03202_ _03620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06565__B _02178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07426_ _02711_ _02918_ _02936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_11_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07240__I _02805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09779__A1 _04496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07357_ _02885_ _00079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06137__S0 _01752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06308_ _01778_ _01923_ _01782_ _01924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08451__A1 _03604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07254__A2 _02807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07288_ _02746_ _02833_ _02836_ _00059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09027_ _03913_ _03959_ _03966_ _00668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06239_ u_cpu.rf_ram.memory\[28\]\[1\] u_cpu.rf_ram.memory\[29\]\[1\] u_cpu.rf_ram.memory\[30\]\[1\]
+ u_cpu.rf_ram.memory\[31\]\[1\] _01631_ _01634_ _01855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06852__I2 u_cpu.rf_ram.memory\[62\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09167__I _03893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11736__CLK net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08203__A1 u_cpu.rf_ram.memory\[19\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10010__A1 _04500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08754__A2 _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06765__A1 _01725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10561__A2 _05088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09929_ _04397_ _04627_ _04633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_93_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09703__A1 _04425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11886__CLK net458 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11822_ _00518_ net477 u_cpu.rf_ram.memory\[143\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07317__I0 u_cpu.rf_ram_if.wdata0_r\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10077__A1 _04561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11753_ _00449_ net481 u_cpu.rf_ram.memory\[142\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10776__I _05219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10704_ u_cpu.rf_ram.memory\[104\]\[0\] _05177_ _05178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11684_ _00388_ net300 u_cpu.rf_ram.memory\[57\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07493__A2 _02970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10635_ _05131_ _05133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_126_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10624__I0 u_arbiter.i_wb_cpu_rdt\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08442__A1 _03598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10566_ _05053_ _05085_ _05092_ _01082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07245__A2 _02806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12305_ _00985_ net502 u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xu_scanchain_local.scan_flop\[40\] u_scanchain_local.module_data_in\[39\] net552 u_arbiter.o_wb_cpu_adr\[2\]
+ net20 u_scanchain_local.module_data_in\[40\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
X_10497_ u_cpu.rf_ram.memory\[97\]\[3\] _05047_ _05050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12236_ _00919_ net264 u_cpu.cpu.immdec.imm19_12_20\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12661__CLK net159 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10001__A1 _01443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12167_ _00850_ net389 u_arbiter.i_wb_cpu_dbus_dat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06300__S0 _01762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06756__A1 _01590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11118_ u_cpu.cpu.genblk3.csr.mstatus_mie _05415_ _05440_ _05441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_1_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12098_ _00781_ net405 u_cpu.rf_ram.memory\[121\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout197_I net202 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11049_ _05347_ _05392_ _05394_ _01263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_42_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10304__A2 _04915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout364_I net365 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07181__A1 _02733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06590_ u_cpu.rf_ram.memory\[56\]\[4\] u_cpu.rf_ram.memory\[57\]\[4\] u_cpu.rf_ram.memory\[58\]\[4\]
+ u_cpu.rf_ram.memory\[59\]\[4\] _01871_ _02099_ _02203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_3690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10068__A1 _04721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout531_I net534 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11609__CLK net236 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06385__B _01999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08260_ _03417_ _03473_ _03480_ _00387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08681__A1 _03019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08156__I _03077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07484__A2 _02973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07211_ _02782_ _02784_ _02785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_105_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12191__CLK net498 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08191_ _03438_ _03440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10615__I0 u_arbiter.i_wb_cpu_rdt\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07142_ _02709_ _02724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11759__CLK net479 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06295__I0 u_cpu.rf_ram.memory\[116\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07073_ u_cpu.rf_ram_if.rdata0\[5\] _02665_ _02668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08984__A2 _03938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06024_ _01575_ _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_47_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08736__A2 _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06747__A1 _01958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10543__A2 _05076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07975_ _03257_ _03299_ _03302_ _00280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09714_ u_arbiter.i_wb_cpu_rdt\[14\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[14\]
+ _04413_ _04439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06926_ u_cpu.cpu.immdec.imm11_7\[0\] _02535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_5_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09161__A2 _04049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09645_ u_arbiter.i_wb_cpu_dbus_dat\[31\] _04380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06857_ u_cpu.rf_ram.memory\[40\]\[7\] u_cpu.rf_ram.memory\[41\]\[7\] u_cpu.rf_ram.memory\[42\]\[7\]
+ u_cpu.rf_ram.memory\[43\]\[7\] _01736_ _02103_ _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_56_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05808_ _01445_ _01449_ _01454_ u_arbiter.o_wb_cpu_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09576_ u_arbiter.i_wb_cpu_dbus_dat\[9\] _04329_ _04333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06788_ _02392_ _02394_ _02396_ _02398_ _01606_ _02399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05722__A2 _01371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10059__A1 _04509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08527_ u_cpu.rf_ram.memory\[72\]\[5\] _03647_ _03651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05739_ u_cpu.cpu.immdec.imm24_20\[0\] _01389_ _01390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_19_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12534__CLK net276 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08458_ u_cpu.rf_ram.memory\[141\]\[0\] _03610_ _03611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08672__A1 u_cpu.rf_ram.memory\[39\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07409_ u_cpu.rf_ram.memory\[78\]\[0\] _02926_ _02927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08389_ _03564_ u_cpu.rf_ram.memory\[9\]\[1\] _03562_ _03565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_13_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10606__I0 u_arbiter.i_wb_cpu_rdt\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10420_ _04990_ _01038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07227__A2 _02796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12684__CLK net232 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10351_ _04948_ _01011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08975__A2 _03935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06986__A1 u_cpu.cpu.branch_op vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10782__A2 _05220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06314__I _01632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10282_ _04906_ _04907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12021_ _00704_ net481 u_cpu.cpu.state.o_cnt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08727__A2 _03767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06738__A1 _02060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10534__A2 _05073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07346__S _02879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10280__B net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout560 net563 net560 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12064__CLK net289 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10298__A1 _01463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10298__B2 u_cpu.cpu.ctrl.o_ibus_adr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06910__A1 _01830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11805_ _00501_ net347 u_cpu.rf_ram.memory\[71\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11736_ _00440_ net149 u_cpu.rf_ram.memory\[15\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08663__A1 u_cpu.rf_ram.memory\[39\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10470__A1 _04419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11667_ _00371_ net114 u_cpu.rf_ram.memory\[5\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10618_ _05122_ _01104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11598_ _00302_ net251 u_cpu.rf_ram.memory\[66\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06277__I0 u_cpu.rf_ram.memory\[104\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08966__A2 _03926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout112_I net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10549_ u_cpu.rf_ram.memory\[95\]\[7\] _05071_ _05082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06977__A1 _02559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11130__I _02745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10773__A2 _05220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09963__C _04662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09915__A1 _04436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09915__B2 _04608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12219_ _00902_ net318 u_cpu.rf_ram.memory\[114\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10525__A2 _05064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12407__CLK net500 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout481_I net483 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07760_ u_cpu.rf_ram.memory\[17\]\[6\] _03158_ _03163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06711_ u_cpu.rf_ram.memory\[92\]\[5\] u_cpu.rf_ram.memory\[93\]\[5\] u_cpu.rf_ram.memory\[94\]\[5\]
+ u_cpu.rf_ram.memory\[95\]\[5\] _02142_ _01915_ _02323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_49_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07691_ _01437_ _03113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_53_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11431__CLK net368 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12557__CLK net212 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09430_ _04225_ _04227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_64_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06642_ _02235_ _02254_ _01810_ _02255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06901__A1 _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09361_ u_cpu.rf_ram.memory\[121\]\[7\] _04172_ _04183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06827__C _01405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[1\]_SE net552 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06573_ _01597_ _02185_ _01795_ _02186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08312_ _03494_ _03513_ _03518_ _00401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_90_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09292_ _04072_ _04130_ _04138_ _00762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07457__A2 _02954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10056__A4 _04736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout25_I net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11581__CLK net339 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10461__A1 _04492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08243_ u_cpu.rf_ram.memory\[58\]\[6\] _03465_ _03470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06760__S0 _01747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07209__A2 _02710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08174_ u_cpu.rf_ram.memory\[60\]\[1\] _03428_ _03430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07125_ _02672_ _02707_ _02671_ u_arbiter.i_wb_cpu_dbus_sel\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08957__A2 _03923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06968__A1 _01411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06968__B2 _02575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10764__A2 _05207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07056_ _02647_ _02656_ _02657_ _00018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06134__I _01609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06007_ _01623_ _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[14\]_SI u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07958_ _03292_ _00273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05943__A2 _01557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09381__S _04185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06909_ u_cpu.rf_ram.memory\[140\]\[7\] u_cpu.rf_ram.memory\[141\]\[7\] u_cpu.rf_ram.memory\[142\]\[7\]
+ u_cpu.rf_ram.memory\[143\]\[7\] _02169_ _01816_ _02519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_28_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07145__A1 _02726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07889_ u_cpu.rf_ram.memory\[74\]\[3\] _03245_ _03247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06579__S0 _02084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09628_ u_arbiter.i_wb_cpu_dbus_dat\[24\] _04295_ _04319_ u_arbiter.i_wb_cpu_dbus_dat\[25\]
+ _04369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_28_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09180__I _03906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09559_ u_arbiter.i_wb_cpu_dbus_dat\[5\] _04289_ _04317_ _04319_ _04320_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_62_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12570_ _01249_ net205 u_cpu.rf_ram.memory\[86\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08645__A1 u_cpu.rf_ram.memory\[138\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06309__I _01426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09693__I0 u_arbiter.i_wb_cpu_rdt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10452__A1 _04468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11521_ _00225_ net430 u_cpu.rf_ram.memory\[129\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10452__B2 _04680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06751__S0 _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11452_ _00156_ net335 u_cpu.rf_ram.memory\[48\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10403_ _04200_ u_cpu.rf_ram.memory\[3\]\[7\] _04972_ _04981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09070__A1 _03977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11383_ _00087_ net215 u_cpu.rf_ram.memory\[80\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06959__A1 _02562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10755__A2 _05207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10334_ u_cpu.cpu.ctrl.o_ibus_adr\[20\] _04936_ _04938_ u_cpu.cpu.ctrl.o_ibus_adr\[21\]
+ _04939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07081__B1 _01411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10265_ u_cpu.rf_ram.memory\[30\]\[1\] _04895_ _04897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10507__A2 _05042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12004_ _00687_ net408 u_cpu.rf_ram.memory\[37\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10196_ u_arbiter.i_wb_cpu_dbus_adr\[8\] u_arbiter.i_wb_cpu_dbus_adr\[7\] _04855_
+ _04856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06026__I3 u_cpu.rf_ram.memory\[27\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11454__CLK net334 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11180__A2 _05481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout390 net391 net390 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_93_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09125__A2 _02563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07439__A2 _02946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10443__A1 _02674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06498__I0 u_cpu.rf_ram.memory\[32\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11719_ _00423_ net332 u_cpu.rf_ram.memory\[52\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout327_I net328 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12699_ u_cpu.rf_ram_if.wdata1_r\[3\] net232 u_cpu.rf_ram_if.wdata1_r\[2\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06742__S0 _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08939__A2 _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09061__A1 _03018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10746__A2 _05201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07611__A2 _03047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08930_ u_cpu.rf_ram.memory\[128\]\[2\] _03904_ _03905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09364__A2 _03166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08861_ _03813_ _03859_ _03861_ _00607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11171__A2 _05466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07812_ _03197_ _03184_ _03198_ _00221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08792_ _03815_ _03817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_111_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11947__CLK net444 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07743_ _03087_ _03143_ _03152_ _00198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_42_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07127__A1 u_cpu.rf_ram_if.genblk1.wtrig0_r vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07674_ _03103_ _00178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09413_ _04145_ _04213_ _04216_ _00805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06625_ u_cpu.rf_ram.memory\[88\]\[4\] u_cpu.rf_ram.memory\[89\]\[4\] u_cpu.rf_ram.memory\[90\]\[4\]
+ u_cpu.rf_ram.memory\[91\]\[4\] _02029_ _01742_ _02238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_77_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06556_ u_cpu.rf_ram.memory\[140\]\[3\] u_cpu.rf_ram.memory\[141\]\[3\] u_cpu.rf_ram.memory\[142\]\[3\]
+ u_cpu.rf_ram.memory\[143\]\[3\] _02169_ _01821_ _02170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09344_ _04172_ _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06129__I _01702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09675__I0 u_arbiter.i_wb_cpu_rdt\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09868__C _04582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10434__A1 _04821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09275_ _02785_ _03970_ _04128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06487_ _02098_ _02100_ _01873_ _02101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06573__B _01795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05968__I _01584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06733__S0 _02169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10985__A2 _05349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11327__CLK net170 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08226_ _03459_ _00374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07850__A2 _03220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05861__A1 _01473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08157_ u_cpu.rf_ram.memory\[61\]\[4\] _03413_ _03418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07108_ _02692_ _02638_ _02696_ _00024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08088_ _03342_ _03369_ _03374_ _00321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07602__A2 _03048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06256__I3 u_cpu.rf_ram.memory\[59\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11477__CLK net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07039_ _02579_ _02642_ _02644_ _02645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10050_ u_cpu.cpu.immdec.imm19_12_20\[2\] _04636_ _04737_ _04742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09355__A2 _04177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07366__A1 _02731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11162__A2 _05469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07118__A1 _02633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10952_ _05332_ _01228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08866__A1 _03821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07669__A2 _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10673__A1 _05142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12102__CLK net444 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10883_ u_cpu.rf_ram.memory\[69\]\[1\] _05290_ _05292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12622_ _01301_ net53 u_cpu.rf_ram.memory\[26\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08618__A1 u_cpu.rf_ram.memory\[143\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06039__I _01595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12553_ _01232_ net212 u_cpu.rf_ram.memory\[85\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09291__A1 u_cpu.rf_ram.memory\[117\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08094__A2 _03370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06724__S0 _01934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09830__A3 _04491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10976__A2 _05337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11504_ _00208_ net295 u_cpu.rf_ram.memory\[40\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12252__CLK net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08254__I _03472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07841__A2 _03217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12484_ _01163_ net40 u_cpu.rf_ram.memory\[105\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11435_ _00139_ net334 u_cpu.rf_ram.memory\[41\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09594__A2 _04338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11366_ _00070_ net122 u_cpu.rf_ram.memory\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10317_ _04928_ _00997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11297_ _05546_ _05551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_79_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09346__A2 _04174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10248_ u_cpu.cpu.bufreg.i_sh_signed _02705_ _02691_ _04884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10179_ u_cpu.rf_ram.memory\[31\]\[7\] _04835_ _04846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[69\]_CLK net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07109__A1 _01431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout277_I net280 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06580__A2 _02192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08429__I _03589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08857__A1 _02722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06707__I1 u_cpu.rf_ram.memory\[117\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10664__A1 _05130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout444_I net447 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06410_ _01423_ _02013_ _02024_ _02025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_50_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07390_ u_cpu.rf_ram.memory\[80\]\[5\] _02901_ _02911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06341_ u_cpu.rf_ram.memory\[12\]\[2\] u_cpu.rf_ram.memory\[13\]\[2\] u_cpu.rf_ram.memory\[14\]\[2\]
+ u_cpu.rf_ram.memory\[15\]\[2\] _01583_ _01841_ _01956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_17_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08085__A2 _03369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06715__S0 _01651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10967__A2 _05340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06096__A1 _01647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09060_ _03988_ _03973_ _03989_ _00678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06272_ _01862_ _01875_ _01887_ _01888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_124_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07832__A2 _03208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06486__I3 u_cpu.rf_ram.memory\[59\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08011_ _03323_ _03324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05843__A1 _01473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11216__I0 _02854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09034__A1 _03033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10719__A2 _05175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09585__A2 _04334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06643__I0 u_cpu.rf_ram.memory\[136\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09962_ _04545_ _04563_ _04660_ _04661_ _04662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__05737__B _01387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09337__A2 _04165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08913_ _03830_ _03883_ _03891_ _00629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_63_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09893_ u_arbiter.i_wb_cpu_rdt\[26\] u_arbiter.i_wb_cpu_rdt\[10\] _01441_ _04599_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11144__A2 _05452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08844_ _03846_ _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10352__B1 _04945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10869__I _04826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05987_ _01597_ _01600_ _01603_ _01604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08775_ _03801_ _03806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12125__CLK net406 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06571__A2 _02183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07726_ _03141_ _03143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08848__A1 _03824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07657_ _03068_ _03090_ _03093_ _00171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07520__A1 _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06608_ u_cpu.rf_ram.memory\[100\]\[4\] u_cpu.rf_ram.memory\[101\]\[4\] u_cpu.rf_ram.memory\[102\]\[4\]
+ u_cpu.rf_ram.memory\[103\]\[4\] _02122_ _01895_ _02221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12275__CLK net533 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07588_ _02996_ _03037_ _03044_ _00151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_70_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09327_ _04140_ _04161_ _04163_ _00772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06539_ _01627_ _02153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11080__A1 _05361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09258_ u_cpu.rf_ram.memory\[34\]\[0\] _04118_ _04119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07823__A2 _03205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05834__A1 u_cpu.cpu.ctrl.o_ibus_adr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08209_ _02786_ _02850_ _03450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__09025__A1 _03910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09189_ _03915_ _04072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_5_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11220_ _02860_ u_cpu.rf_ram.memory\[0\]\[3\] _05501_ _05505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09576__A2 _04329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08802__I _03497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06750__C _01807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11151_ _05462_ _05447_ _05463_ _01296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10102_ _04469_ _04783_ _04787_ _04511_ _04788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_68_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11082_ _05363_ _05405_ _05413_ _01277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11135__A2 _05452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10033_ _04402_ _04502_ _04726_ _04509_ _04727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_103_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08000__A2 _03316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10343__B1 _04938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06937__I1 _02545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07354__S _02879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06562__A2 _02175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08249__I _03472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11984_ _00674_ net438 u_cpu.rf_ram.memory\[123\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07153__I _02734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10935_ u_cpu.rf_ram.memory\[59\]\[6\] _05318_ _05323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07511__A1 _02992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10866_ _04823_ _05280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12605_ _01284_ net378 u_cpu.cpu.genblk3.csr.mstatus_mpie vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08067__A2 _03356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09264__A1 _04063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11642__CLK net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10797_ u_cpu.rf_ram.memory\[106\]\[2\] _05236_ _05237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11071__A1 _05352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07102__B _02691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12536_ _01215_ net278 u_cpu.rf_ram.memory\[59\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06468__I3 u_cpu.rf_ram.memory\[19\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05825__A1 u_cpu.cpu.ctrl.o_ibus_adr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09016__A1 _03894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12467_ _01146_ net45 u_cpu.rf_ram.memory\[99\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09808__I _04527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11792__CLK net373 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11418_ _00122_ net291 u_cpu.rf_ram.memory\[44\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12398_ _01077_ net44 u_cpu.rf_ram.memory\[96\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06625__I0 u_cpu.rf_ram.memory\[88\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11349_ _00053_ net69 u_cpu.rf_ram.memory\[18\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09319__A2 _04143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout394_I net395 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05910_ u_arbiter.i_wb_cpu_dbus_adr\[23\] _01512_ _01536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06890_ _01740_ _02499_ _01744_ _02500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10334__B1 _04938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05841_ _01452_ _01481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_fanout561_I net562 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07750__A1 _03068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08560_ u_cpu.rf_ram.memory\[71\]\[1\] _03669_ _03672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08159__I _03080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05772_ _01422_ _01423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_66_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07063__I _01401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10637__A1 _05130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07511_ _02992_ _02984_ _02993_ _00125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_63_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08491_ u_cpu.rf_ram.memory\[140\]\[6\] _03625_ _03630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06305__A2 _01920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07442_ _02904_ _02942_ _02948_ _00101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout18 net19 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_62_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout29 net31 net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XFILLER_50_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07373_ u_cpu.rf_ram.memory\[80\]\[1\] _02894_ _02898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08058__A2 _02923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09255__A1 _02722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11062__A1 _05363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09112_ _03980_ _04015_ _04021_ _00698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06324_ _01760_ _01926_ _01939_ _01940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__06164__S1 _01780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09043_ _03971_ _03978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09007__A1 _03913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06255_ _01673_ _01871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_102_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06851__B _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06186_ _01706_ _01803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_11_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07569__A1 u_cpu.rf_ram.memory\[41\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08230__A2 _03462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10092__C _04575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07238__I _02803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09945_ _04469_ _04638_ _04646_ _04466_ _04647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_132_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11117__A2 _02567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06792__A2 _02402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09876_ u_cpu.rf_ram.memory\[114\]\[0\] _04589_ _04590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05981__I _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11515__CLK net321 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09730__A2 _04454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08827_ u_cpu.rf_ram.memory\[132\]\[3\] _03839_ _03841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07741__A1 _03084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08758_ u_cpu.rf_ram.memory\[135\]\[3\] _03794_ _03796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07709_ _03121_ _03129_ _03130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08297__A2 _03495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08689_ _03493_ _03752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11665__CLK net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06147__I2 u_cpu.rf_ram.memory\[94\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10720_ _05148_ _05177_ _05186_ _01142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09246__A1 _04066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10651_ _04826_ _05144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09797__A2 _04418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10582_ u_cpu.rf_ram.memory\[28\]\[1\] _05101_ _05103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05807__A1 u_arbiter.i_wb_cpu_dbus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12321_ _01001_ net532 u_cpu.cpu.ctrl.o_ibus_adr\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10800__A1 _05209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06480__A1 _01656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12252_ _00935_ net93 u_cpu.rf_ram.memory\[31\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11203_ _05454_ _05489_ _05495_ _01316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_12183_ _00866_ net389 u_arbiter.i_wb_cpu_dbus_dat\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11098__C _02684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11134_ _05445_ _05452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_7_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07980__A1 _03262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06783__A2 _02393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11065_ _05300_ _03166_ _05403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09363__I _02845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10016_ _04680_ _04452_ _04710_ _04612_ _04711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_76_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10867__A1 u_cpu.rf_ram.memory\[108\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06535__A2 _02148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05969__S1 _01585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06091__S0 _01705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09485__A1 _04244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11967_ _00663_ net464 u_cpu.rf_ram.memory\[124\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10918_ _05286_ _05303_ _05312_ _01214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11898_ _00594_ net471 u_cpu.rf_ram.memory\[132\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06394__S1 _01895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout142_I net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10849_ _05217_ _05258_ _05267_ _01190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11133__I _02751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11044__A1 _05365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[40\]_SE net552 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07799__A1 u_cpu.rf_ram.memory\[119\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12519_ _01198_ net171 u_cpu.rf_ram.memory\[108\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout407_I net413 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08460__A2 _03610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06040_ _01620_ _01657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_132_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06861__I3 u_cpu.rf_ram.memory\[39\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.output_buffers\[2\] u_scanchain_local.data_out_i u_scanchain_local.data_out
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11538__CLK net234 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout208 net209 net208 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__09960__A2 _04659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout219 net223 net219 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_114_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07991_ _03311_ _03312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06774__A2 _02384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09730_ _04403_ _04454_ _04455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06942_ _02534_ _02548_ _02550_ _02551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10413__S _04983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10858__A1 _05273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09661_ _04247_ _04384_ _04390_ _00879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06873_ _01802_ _02482_ _02483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08612_ u_cpu.rf_ram.memory\[143\]\[3\] _03704_ _03706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05824_ _01463_ _01464_ u_cpu.cpu.ctrl.o_ibus_adr\[6\] _01467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09592_ u_arbiter.i_wb_cpu_rdt\[12\] _04334_ _04344_ u_arbiter.i_wb_cpu_dbus_dat\[12\]
+ _04345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_97_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout55_I net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08543_ u_cpu.rf_ram.memory\[73\]\[3\] _03659_ _03661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05755_ _01404_ _01405_ _01406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_97_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09476__A1 _02830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06909__S0 _02169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06846__B _01588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11283__A1 _02906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08474_ _03606_ _03610_ _03619_ _00462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07521__I _02915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07425_ _02916_ _02926_ _02935_ _00097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09228__A1 _04068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07356_ _02867_ u_cpu.rf_ram.memory\[7\]\[5\] _02878_ _02885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_17_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06307_ u_cpu.rf_ram.memory\[84\]\[1\] u_cpu.rf_ram.memory\[85\]\[1\] u_cpu.rf_ram.memory\[86\]\[1\]
+ u_cpu.rf_ram.memory\[87\]\[1\] _01922_ _01780_ _01923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_40_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07287_ u_cpu.rf_ram.memory\[20\]\[1\] _02834_ _02836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08451__A2 _03591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09448__I _03893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06462__A1 _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09026_ u_cpu.rf_ram.memory\[124\]\[5\] _03962_ _03966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06238_ _01619_ _01853_ _01628_ _01854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_105_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06852__I3 u_cpu.rf_ram.memory\[63\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06169_ _01683_ _01786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_65_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10397__I0 _04194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09384__S _04185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12463__CLK net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09928_ _04629_ _04631_ _04632_ _04557_ _00904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_28_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09183__I _03909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09703__A2 _04426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10849__A1 _05217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09859_ u_arbiter.i_wb_cpu_rdt\[22\] u_arbiter.i_wb_cpu_rdt\[6\] _01446_ _04574_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_8_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07714__A1 _03119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11821_ _00517_ net486 u_cpu.rf_ram.memory\[143\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07317__I1 u_cpu.rf_ram_if.wdata1_r\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10077__A2 _04502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11274__A1 _02888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11752_ _00448_ net479 u_cpu.rf_ram.memory\[142\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[63\]_SE net556 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06376__S1 _01699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06475__C _01428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10703_ _05175_ _05177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_14_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09219__A1 _04056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11683_ _00387_ net324 u_cpu.rf_ram.memory\[57\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10634_ _05131_ _05132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10624__I1 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08442__A2 _03590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10565_ u_cpu.rf_ram.memory\[96\]\[5\] _05088_ _05092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12304_ _00984_ net500 u_arbiter.i_wb_cpu_ibus_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06453__A1 _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10496_ _04820_ _05049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[33\] u_arbiter.i_wb_cpu_rdt\[30\] net550 u_arbiter.i_wb_cpu_dbus_dat\[27\]
+ net17 u_arbiter.i_wb_cpu_rdt\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
X_12235_ _00918_ net263 u_cpu.cpu.immdec.imm19_12_20\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10001__A2 u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12166_ _00849_ net391 u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06756__A2 _02366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06300__S1 _01915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11117_ _04952_ _02567_ _05440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_12097_ _00780_ net410 u_cpu.rf_ram.memory\[121\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11048_ u_cpu.rf_ram.memory\[87\]\[0\] _05393_ _05394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08638__S _03711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11980__CLK net254 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07181__A2 _02758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout357_I net366 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08505__I0 _03570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11265__A1 _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08437__I _03589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08130__A1 u_cpu.rf_ram.memory\[62\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout524_I net527 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12336__CLK net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08681__A2 _03698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07210_ _02783_ _02715_ _02784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__11017__A1 u_cpu.rf_ram.memory\[86\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08190_ _03438_ _03439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06819__I0 u_cpu.rf_ram.memory\[136\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07141_ _02722_ _02723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_88_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11360__CLK net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07072_ _01430_ _02654_ _02667_ _00011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06295__I1 u_cpu.rf_ram.memory\[117\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12486__CLK net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06023_ _01639_ _01640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08197__A1 u_cpu.rf_ram.memory\[19\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05745__B _01388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07974_ u_cpu.rf_ram.memory\[68\]\[1\] _03300_ _03302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09713_ _04437_ _04418_ _04438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06925_ u_cpu.cpu.alu.i_rs1 u_cpu.cpu.alu.add_cy_r _02534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09644_ _04376_ _04322_ _04329_ _04378_ _04379_ _00873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_67_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06856_ _02459_ _02461_ _02463_ _02465_ _01427_ _02466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_82_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05807_ u_arbiter.i_wb_cpu_dbus_adr\[2\] _01453_ _01454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09575_ _04330_ _04332_ _00851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09449__A1 _03002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06787_ _01720_ _02397_ _01663_ _02398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05722__A3 _01372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10059__A2 _04548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08526_ _03600_ _03643_ _03650_ _00483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11256__A1 _02896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05738_ _01368_ _01378_ _01388_ _01389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_51_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08457_ _03608_ _03610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_24_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11008__A1 u_cpu.rf_ram.memory\[86\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07408_ _02924_ _02926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08388_ _02854_ _03564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_17_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07339_ _02873_ u_cpu.rf_ram.memory\[1\]\[7\] _02851_ _02874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06286__I1 u_cpu.rf_ram.memory\[125\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10350_ _01547_ _04943_ _04945_ u_cpu.cpu.ctrl.o_ibus_adr\[28\] _04948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_139_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06986__A2 u_cpu.cpu.decode.opcode\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09009_ _03916_ _03947_ _03955_ _00661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10281_ _04905_ _04906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11853__CLK net510 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08188__A1 _03423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12020_ _00703_ net379 u_cpu.cpu.state.stage_two_req vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06738__A2 _02349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout550 net551 net550 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__12209__CLK net373 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout561 net562 net561 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10298__A2 _04915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08360__A1 _03507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06597__S1 _02109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06910__A2 _02519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11804_ _00500_ net348 u_cpu.rf_ram.memory\[71\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11247__A1 _05460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08112__A1 u_cpu.rf_ram.memory\[63\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_37_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11735_ _00439_ net136 u_cpu.rf_ram.memory\[15\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10470__A2 _04452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11666_ _00370_ net70 u_cpu.rf_ram.memory\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10617_ u_arbiter.i_wb_cpu_rdt\[25\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[9\]
+ _05117_ _05122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11597_ _00301_ net251 u_cpu.rf_ram.memory\[66\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10548_ _05055_ _05073_ _05081_ _01075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout105_I net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10479_ _04493_ _04491_ _05035_ _05036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_142_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12218_ _00901_ net316 u_cpu.rf_ram.memory\[114\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09915__A2 _04566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07926__A1 _03270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06729__A2 _02331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12149_ _00832_ net317 u_cpu.rf_ram.memory\[116\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06710_ _01647_ _02312_ _02321_ _02322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_49_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06037__S0 _01651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07690_ _03111_ _03112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_77_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06641_ _02026_ _02244_ _02253_ _02254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_65_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11238__A1 u_cpu.rf_ram.memory\[98\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09360_ _04156_ _04174_ _04182_ _00786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06572_ u_cpu.rf_ram.memory\[0\]\[4\] u_cpu.rf_ram.memory\[1\]\[4\] u_cpu.rf_ram.memory\[2\]\[4\]
+ u_cpu.rf_ram.memory\[3\]\[4\] _02074_ _01585_ _02185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_17_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11726__CLK net416 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08311_ u_cpu.rf_ram.memory\[55\]\[2\] _03517_ _03518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09291_ u_cpu.rf_ram.memory\[117\]\[6\] _04133_ _04138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09851__A1 _04432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08654__A2 _03726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08242_ _03419_ _03462_ _03469_ _00380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout18_I net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06760__S1 _01748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11876__CLK net516 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08173_ _03405_ _03427_ _03429_ _00351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06417__A1 _01766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07124_ _01369_ _02672_ _02671_ u_arbiter.i_wb_cpu_dbus_sel\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06512__S1 _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07055_ _02646_ u_cpu.rf_ram_if.rdata1\[4\] _02657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_12_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06006_ u_cpu.raddr\[1\] _01623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07917__A1 _03264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08590__A1 _03673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07246__I _02805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06150__I _01704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07957_ _02858_ u_cpu.rf_ram.memory\[6\]\[2\] _03289_ _03292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12501__CLK net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06908_ _01825_ _02517_ _02518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_28_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07888_ _03188_ _03241_ _03246_ _00249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09461__I _03906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08342__A1 _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06579__S1 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09627_ u_arbiter.i_wb_cpu_rdt\[24\] _04312_ _04368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06839_ u_cpu.rf_ram.memory\[20\]\[7\] u_cpu.rf_ram.memory\[21\]\[7\] u_cpu.rf_ram.memory\[22\]\[7\]
+ u_cpu.rf_ram.memory\[23\]\[7\] _01631_ _01634_ _02449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_56_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09558_ _04318_ _04319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_58_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12651__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08509_ _03574_ u_cpu.rf_ram.memory\[13\]\[6\] _03632_ _03640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_19_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09489_ _04249_ _04258_ _04265_ _00832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_12_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11520_ _00224_ net430 u_cpu.rf_ram.memory\[129\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10452__A2 _04510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08805__I _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06751__S1 _01965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11451_ _00155_ net333 u_cpu.rf_ram.memory\[48\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10402_ _04980_ _01030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11382_ _00086_ net185 u_cpu.rf_ram.memory\[80\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06959__A2 _02563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07081__A1 _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10333_ _04908_ _04938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_106_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10264_ _04808_ _04894_ _04896_ _00976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12003_ _00686_ net415 u_cpu.rf_ram.memory\[38\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10195_ _04848_ _04855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_78_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08581__A1 _03272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12181__CLK net389 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout380 net381 net380 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_43_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06592__B1 _02202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout391 net392 net391 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_4_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09371__I _02857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11749__CLK net256 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10140__A1 _04817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10691__A2 _05168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11899__CLK net471 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09833__A1 _04548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10443__A2 _02704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06498__I1 u_cpu.rf_ram.memory\[33\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11718_ _00422_ net415 u_cpu.rf_ram.memory\[53\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12698_ u_cpu.rf_ram_if.wdata1_r\[2\] net140 u_cpu.rf_ram_if.wdata1_r\[1\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06742__S1 _01592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout222_I net223 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11649_ _00353_ net215 u_cpu.rf_ram.memory\[60\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09061__A2 _03286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07072__A1 _01430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08860_ u_cpu.rf_ram.memory\[130\]\[0\] _03860_ _03861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07811_ u_cpu.rf_ram.memory\[119\]\[6\] _03189_ _03198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08791_ _03815_ _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10421__S _04982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07742_ u_cpu.rf_ram.memory\[16\]\[7\] _03141_ _03152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07127__A2 _01387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09372__I0 _04190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12674__CLK net256 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06838__C _01807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07673_ _02846_ u_cpu.rf_ram.memory\[4\]\[0\] _03102_ _03103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10131__A1 _04808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08875__A2 _03858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09412_ u_cpu.rf_ram.memory\[112\]\[1\] _04214_ _04216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06430__S0 _01934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06624_ _01761_ _02236_ _02237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06886__A1 _01647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09343_ _03019_ _03970_ _04172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06555_ _01813_ _02169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_52_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09824__A1 _04516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09274_ _04074_ _04118_ _04127_ _00755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10434__A2 _04993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06486_ u_cpu.rf_ram.memory\[56\]\[3\] u_cpu.rf_ram.memory\[57\]\[3\] u_cpu.rf_ram.memory\[58\]\[3\]
+ u_cpu.rf_ram.memory\[59\]\[3\] _01871_ _02099_ _02100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06733__S1 _01816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08225_ _02873_ u_cpu.rf_ram.memory\[5\]\[7\] _03450_ _03459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_53_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09588__B1 _04331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06145__I _01612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08156_ _03077_ _03417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07107_ _02528_ _02695_ _02696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08087_ u_cpu.rf_ram.memory\[29\]\[2\] _03373_ _03374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07038_ _02613_ _02603_ _02643_ _02578_ _02644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_115_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07366__A2 _02891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10370__A1 u_cpu.rf_ram.memory\[109\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08989_ _03916_ _03935_ _03943_ _00653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07118__A2 _02703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10951_ _04196_ u_cpu.rf_ram.memory\[10\]\[5\] _05325_ _05332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06177__I0 u_cpu.rf_ram.memory\[68\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10122__A1 _04026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08866__A2 _03859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10673__A2 _05151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06421__S0 _01922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10882_ _05268_ _05289_ _05291_ _01199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12621_ _01300_ net51 u_cpu.rf_ram.memory\[26\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09815__A1 _04505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08618__A2 _03704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09140__B _02699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12552_ _01231_ net212 u_cpu.rf_ram.memory\[85\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07677__I0 _02858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06724__S1 _01763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11503_ _00207_ net295 u_cpu.rf_ram.memory\[40\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12483_ _01162_ net40 u_cpu.rf_ram.memory\[105\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06055__I _01671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11434_ _00138_ net327 u_cpu.rf_ram.memory\[41\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12547__CLK net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11421__CLK net297 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11365_ _00069_ net121 u_cpu.rf_ram.memory\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10316_ u_cpu.cpu.ctrl.o_ibus_adr\[13\] _04922_ _04924_ _01502_ _04928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_106_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11296_ _02896_ _05547_ _05550_ _01354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10247_ _04882_ _02691_ _04883_ _00972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08554__A1 _02876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11571__CLK net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12697__CLK net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10361__A1 _02545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10178_ _04830_ _04837_ _04845_ _00941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10241__S _04848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06660__S0 _02074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07614__I _03059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10113__A1 _04511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout172_I net173 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08857__A2 _03814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06707__I2 u_cpu.rf_ram.memory\[118\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06412__S0 _01762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10664__A2 _05151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_fanout437_I net442 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06340_ _01570_ _01954_ _01955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12077__CLK net310 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06715__S1 _02033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06271_ _01878_ _01881_ _01884_ _01886_ _01711_ _01887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__06096__A2 _01682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07293__A1 _02758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08010_ _02723_ _02923_ _03323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09034__A2 _03970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06479__S0 _01657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07596__A2 _03049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09961_ _04528_ _04567_ _04615_ _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_48_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08912_ u_cpu.rf_ram.memory\[22\]\[6\] _03886_ _03891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09892_ _04255_ _04589_ _04598_ _00902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout85_I net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08545__A1 u_cpu.rf_ram.memory\[73\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08843_ _03819_ _03847_ _03850_ _00600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08774_ _03750_ _03802_ _03805_ _00576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05986_ _01602_ _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07725_ _03141_ _03142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08848__A2 _03847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06403__S0 _01741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10655__A2 _05138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07656_ u_cpu.rf_ram.memory\[50\]\[1\] _03091_ _03093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07520__A2 _02985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06607_ _02004_ _02219_ _01723_ _02220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_90_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07587_ u_cpu.rf_ram.memory\[43\]\[5\] _03040_ _03044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05979__I _01595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09326_ u_cpu.rf_ram.memory\[118\]\[0\] _04162_ _04163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06538_ u_cpu.rf_ram.memory\[84\]\[3\] u_cpu.rf_ram.memory\[85\]\[3\] u_cpu.rf_ram.memory\[86\]\[3\]
+ u_cpu.rf_ram.memory\[87\]\[3\] _01922_ _02151_ _02152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_55_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09257_ _04116_ _04118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11444__CLK net326 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06469_ _02081_ _02082_ _01970_ _02083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_120_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09387__S _04185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08208_ _03423_ _03440_ _03449_ _00366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05834__A2 u_cpu.cpu.ctrl.o_ibus_adr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09025__A2 _03958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09188_ _04070_ _04059_ _04071_ _00724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08139_ _03353_ _03395_ _03404_ _00342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09186__I _03912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11594__CLK net246 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07587__A2 _03040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11150_ u_cpu.rf_ram.memory\[27\]\[7\] _05445_ _05463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10101_ _04784_ _04786_ _04699_ _04787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10125__I _02738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11081_ u_cpu.rf_ram.memory\[88\]\[6\] _05408_ _05413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[1\]_D u_cpu.cpu.genblk3.csr.i_mtip vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08536__A1 u_cpu.rf_ram.memory\[73\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10032_ _04721_ _04489_ _04726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10343__A1 _01537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10343__B2 u_cpu.cpu.ctrl.o_ibus_adr\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10894__A2 _05293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11983_ _00673_ net410 u_cpu.rf_ram.memory\[123\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10646__A2 _05138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10934_ _05282_ _05315_ _05322_ _01220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_16_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07511__A2 _02984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10865_ _05278_ _05270_ _05279_ _01194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12604_ _01283_ net378 u_cpu.cpu.genblk3.csr.mcause31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10796_ _05231_ _05236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xu_scanchain_local.scan_flop\[63\] u_scanchain_local.module_data_in\[62\] net556 u_arbiter.o_wb_cpu_adr\[25\]
+ net24 u_scanchain_local.module_data_in\[63\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_13_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12535_ _01214_ net277 u_cpu.rf_ram.memory\[84\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07275__A1 u_cpu.rf_ram.memory\[18\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05825__A2 _01463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12466_ _01145_ net46 u_cpu.rf_ram.memory\[99\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09016__A2 _03958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11417_ _00121_ net225 u_cpu.rf_ram.memory\[45\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12397_ _01076_ net200 u_cpu.rf_ram.memory\[95\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07578__A2 _03037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06625__I1 u_cpu.rf_ram.memory\[89\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11348_ _00052_ net67 u_cpu.rf_ram.memory\[18\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10582__A1 u_cpu.rf_ram.memory\[28\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06881__S0 _02133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11279_ _02899_ _05535_ _05540_ _01347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08527__A1 u_cpu.rf_ram.memory\[72\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout387_I net388 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10185__I1 u_arbiter.i_wb_cpu_dbus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05840_ u_cpu.cpu.ctrl.o_ibus_adr\[9\] _01477_ _01480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_39_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07750__A2 _03154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout554_I net556 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05771_ _01420_ _01421_ _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_81_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05761__A1 _01409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07510_ u_cpu.rf_ram.memory\[44\]\[3\] _02990_ _02993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08490_ _03602_ _03622_ _03629_ _00468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10637__A2 _05132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07441_ u_cpu.rf_ram.memory\[42\]\[3\] _02946_ _02948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11467__CLK net301 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout19 net35 net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_90_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05799__I _01441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07372_ _02896_ _02897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09255__A2 _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09111_ u_cpu.rf_ram.memory\[36\]\[3\] _04019_ _04021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06323_ _01928_ _01933_ _01936_ _01938_ _01807_ _01939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__11062__A2 _05393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09042_ _03902_ _03977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06254_ _01666_ _01869_ _01870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08903__I _03881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09007__A2 _03947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07018__A1 _01374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06185_ _01777_ _01802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09963__B1 _04486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10573__A1 u_arbiter.i_wb_cpu_ack vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09944_ _04582_ _04641_ _04644_ _04645_ _04526_ _04646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_67_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06872__S0 _02122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09734__I _04458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08518__A1 u_cpu.rf_ram.memory\[72\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09875_ _04587_ _04589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_63_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09191__A1 _04072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08826_ _03821_ _03835_ _03840_ _00593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12242__CLK net383 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07741__A2 _03143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08757_ _03752_ _03790_ _03795_ _00569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05752__A1 u_cpu.cpu.immdec.imm24_20\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05969_ u_cpu.rf_ram.memory\[12\]\[0\] u_cpu.rf_ram.memory\[13\]\[0\] u_cpu.rf_ram.memory\[14\]\[0\]
+ u_cpu.rf_ram.memory\[15\]\[0\] _01583_ _01585_ _01586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_2616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07708_ _03124_ _03128_ _03129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08688_ _03750_ _03747_ _03751_ _00544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07639_ _02767_ _03080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10650_ _05142_ _05132_ _05143_ _01115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09246__A2 _04105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09309_ u_cpu.rf_ram.memory\[120\]\[3\] _04148_ _04151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10581_ _05039_ _05100_ _05102_ _01087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12320_ _01000_ net532 u_cpu.cpu.ctrl.o_ibus_adr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05807__A2 _01453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[68\]_CLK net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10800__A2 _05232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12251_ _00934_ net274 u_cpu.rf_ram.memory\[32\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08757__A1 _03752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11202_ u_cpu.rf_ram.memory\[24\]\[3\] _05493_ _05495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09954__B1 _04560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12182_ _00865_ net389 u_arbiter.i_wb_cpu_dbus_dat\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10564__A1 _05051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06768__B1 _02376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11133_ _02751_ _05451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06863__S0 _01767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07980__A2 _03299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11064_ _05365_ _05393_ _05402_ _01270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09182__A1 _04066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10015_ _04709_ _04710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_49_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06615__S0 _01674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10867__A2 _05276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07164__I _02744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07732__A2 _03146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06091__S1 _01707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11966_ _00662_ net453 u_cpu.rf_ram.memory\[125\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09485__A2 _04258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10917_ u_cpu.rf_ram.memory\[84\]\[7\] _05301_ _05312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11897_ _00593_ net470 u_cpu.rf_ram.memory\[132\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[34\]_D u_arbiter.i_wb_cpu_rdt\[31\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06508__I _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10848_ u_cpu.rf_ram.memory\[83\]\[7\] _05256_ _05267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07248__A1 _02752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout135_I net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10779_ u_cpu.rf_ram.memory\[105\]\[3\] _05224_ _05226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06952__B _02557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08996__A1 _03894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12518_ _01197_ net203 u_cpu.rf_ram.memory\[108\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06671__C _01784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12115__CLK net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12449_ _01128_ net88 u_cpu.rf_ram.memory\[103\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout302_I net303 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08748__A1 _02876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06243__I _01587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10555__A1 _05039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06854__S0 _01729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07990_ _03272_ _03310_ _03311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout209 net214 net209 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_119_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12265__CLK net515 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06941_ _02549_ u_cpu.cpu.alu.add_cy_r _02550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09660_ u_cpu.rf_ram.memory\[113\]\[3\] _04388_ _04390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06606__S0 _02005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06872_ u_cpu.rf_ram.memory\[100\]\[7\] u_cpu.rf_ram.memory\[101\]\[7\] u_cpu.rf_ram.memory\[102\]\[7\]
+ u_cpu.rf_ram.memory\[103\]\[7\] _02122_ _01576_ _02482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_28_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10858__A2 _05270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08611_ _03673_ _03700_ _03705_ _00513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05823_ _01456_ _01465_ _01466_ u_arbiter.o_wb_cpu_adr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09591_ _04294_ _04344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06782__I0 u_cpu.rf_ram.memory\[104\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08542_ _03595_ _03655_ _03660_ _00489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05754_ _01378_ _01388_ _01401_ _01405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_70_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout48_I net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09476__A2 _04224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06909__S1 _01816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07487__A1 _02907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08473_ u_cpu.rf_ram.memory\[141\]\[7\] _03608_ _03619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07424_ u_cpu.rf_ram.memory\[78\]\[7\] _02924_ _02935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06418__I _01652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[25\]_D u_arbiter.i_wb_cpu_rdt\[22\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07239__A1 _02731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07355_ _02884_ _00078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11035__A2 _05384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08987__A1 _03913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06306_ _01572_ _01922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_30_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07286_ _02740_ _02833_ _02835_ _00058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09025_ _03910_ _03958_ _03965_ _00667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06462__A2 _02075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06237_ u_cpu.rf_ram.memory\[16\]\[1\] u_cpu.rf_ram.memory\[17\]\[1\] u_cpu.rf_ram.memory\[18\]\[1\]
+ u_cpu.rf_ram.memory\[19\]\[1\] _01852_ _01625_ _01853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_121_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08739__A1 _03755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12608__CLK net360 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06153__I _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06168_ _01765_ _01771_ _01776_ _01783_ _01784_ _01785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_116_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10546__A1 _05053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07411__A1 u_cpu.rf_ram.memory\[78\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10604__S _05111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06845__S0 _01622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06099_ _01638_ _01716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_132_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09464__I _03909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05992__I _01397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09927_ u_cpu.cpu.immdec.imm24_20\[0\] _04628_ _04632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09164__A1 _03986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09858_ _02571_ _04398_ _04573_ _00893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09703__A3 _04427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08911__A1 _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06368__I3 u_cpu.rf_ram.memory\[59\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08809_ u_cpu.rf_ram.memory\[133\]\[5\] _03822_ _03829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09789_ _04481_ _04511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06773__I0 u_cpu.rf_ram.memory\[36\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11820_ _00516_ net485 u_cpu.rf_ram.memory\[143\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08808__I _03503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11751_ _00447_ net479 u_cpu.rf_ram.memory\[142\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07478__A1 _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10702_ _05175_ _05176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10482__B1 _05037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[16\]_D u_arbiter.i_wb_cpu_rdt\[13\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11682_ _00386_ net324 u_cpu.rf_ram.memory\[57\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10633_ _02785_ _04959_ _05131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12138__CLK net403 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08978__A1 _03900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10564_ _05051_ _05084_ _05091_ _01081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12303_ _00023_ net500 u_cpu.cpu.ctrl.pc_plus_4_cy_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06453__A2 _02066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07650__A1 _03087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10495_ _05046_ _05041_ _05048_ _01055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07159__I _02732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12288__CLK net523 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12234_ _00917_ net263 u_cpu.cpu.immdec.imm19_12_20\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10537__A1 _05044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_scanchain_local.scan_flop\[26\] u_arbiter.i_wb_cpu_rdt\[23\] net545 u_arbiter.i_wb_cpu_dbus_dat\[20\]
+ net13 u_arbiter.i_wb_cpu_rdt\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
X_12165_ _00848_ net390 u_arbiter.i_wb_cpu_dbus_dat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06836__S0 _02074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09374__I _02860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11116_ u_cpu.cpu.genblk3.csr.mstatus_mpie _01378_ _01394_ _05439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12096_ _00779_ net408 u_cpu.rf_ram.memory\[118\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09155__A1 u_cpu.rf_ram.memory\[91\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07108__B _02696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11047_ _05391_ _05393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06012__B _01628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08902__A1 _03819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07622__I _02745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09702__I0 u_arbiter.i_wb_cpu_rdt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout252_I net253 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11265__A2 _05524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11949_ _00645_ net461 u_cpu.rf_ram.memory\[127\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06141__B2 _01756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06531__I3 u_cpu.rf_ram.memory\[91\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10983__I _02745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11017__A2 _05372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout517_I net520 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08969__A1 _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07140_ _02716_ _02721_ _02722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06819__I1 u_cpu.rf_ram.memory\[137\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11505__CLK net302 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09993__B _04619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07071_ u_cpu.rf_ram_if.rdata0\[4\] _02665_ _02667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06444__A2 _02058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07641__A1 u_cpu.rf_ram.memory\[47\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06295__I2 u_cpu.rf_ram.memory\[118\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06022_ _01638_ _01639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_127_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10528__A1 _05055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07944__A2 _03278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05745__C _01367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07973_ _03252_ _03299_ _03301_ _00279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09712_ u_arbiter.i_wb_cpu_rdt\[0\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[0\]
+ _01439_ _04437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06924_ u_arbiter.i_wb_cpu_dbus_we u_cpu.cpu.bufreg.i_sh_signed _02531_ _02532_ _02533_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_132_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09697__A2 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09643_ u_arbiter.i_wb_cpu_rdt\[29\] _04300_ _04379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06855_ _02098_ _02464_ _01695_ _02465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10700__A1 _05148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06755__I0 u_cpu.rf_ram.memory\[28\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06904__B1 _02511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05806_ _01452_ _01453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09574_ u_arbiter.i_wb_cpu_rdt\[7\] _04312_ _04331_ u_arbiter.i_wb_cpu_dbus_dat\[7\]
+ _04332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_58_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06786_ u_cpu.rf_ram.memory\[96\]\[6\] u_cpu.rf_ram.memory\[97\]\[6\] u_cpu.rf_ram.memory\[98\]\[6\]
+ u_cpu.rf_ram.memory\[99\]\[6\] _02125_ _01693_ _02397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_93_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09449__A2 _04224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08525_ u_cpu.rf_ram.memory\[72\]\[4\] _03647_ _03650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05737_ _01380_ _01383_ _01387_ _01388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__11256__A2 _05523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08456_ _03608_ _03609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07407_ _02924_ _02925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_17_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11008__A2 _05369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08387_ _03563_ _00431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07338_ _02872_ _02873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12430__CLK net363 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10767__A1 u_cpu.rf_ram.memory\[79\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09621__A2 _04352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07269_ u_cpu.rf_ram.memory\[18\]\[3\] _02822_ _02824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09395__S _04203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09008_ u_cpu.rf_ram.memory\[125\]\[6\] _03950_ _03955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10280_ _02528_ _02705_ net2 _04905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__10519__A1 u_cpu.rf_ram.memory\[94\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08188__A2 _03428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11192__A1 _05098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout540 net5 net540 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout551 net565 net551 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_76_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10133__I _04813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout562 net563 net562 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_8_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[30\]_SE net547 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07699__A1 _02569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06767__B _01695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08360__A2 _03538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11803_ _00499_ net369 u_cpu.rf_ram.memory\[71\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08499__I0 _03564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11247__A2 _05512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08112__A2 _03386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11734_ _00438_ net143 u_cpu.rf_ram.memory\[9\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06058__I _01658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11528__CLK net511 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11665_ _00369_ net58 u_cpu.rf_ram.memory\[5\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10616_ _05121_ _01103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11596_ _00300_ net251 u_cpu.rf_ram.memory\[66\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09612__A2 _04352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10758__A1 u_cpu.rf_ram.memory\[79\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11678__CLK net299 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10547_ u_cpu.rf_ram.memory\[95\]\[6\] _05076_ _05081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10478_ _04567_ _05034_ _04487_ _04575_ _05035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_68_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08179__A2 _03431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12217_ _00900_ net316 u_cpu.rf_ram.memory\[114\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08423__I0 _03574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11183__A1 _05454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07926__A2 _03255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12148_ _00831_ net317 u_cpu.rf_ram.memory\[116\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05937__A1 _01489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10930__A1 _05278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12079_ _00762_ net319 u_cpu.rf_ram.memory\[117\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09832__I _04527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06037__S1 _01653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout467_I net473 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12303__CLK net500 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08351__A2 _03541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06640_ _02246_ _02248_ _02250_ _02252_ _02050_ _02253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_20_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06571_ _01958_ _02183_ _02184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11238__A2 _05515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09300__A1 _04140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08103__A2 _03383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08310_ _03512_ _03517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09290_ _04070_ _04130_ _04137_ _00761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12453__CLK net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09851__A2 _04477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08241_ u_cpu.rf_ram.memory\[58\]\[5\] _03465_ _03469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10419__S _04982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08172_ u_cpu.rf_ram.memory\[60\]\[0\] _03428_ _03429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10749__A1 _05204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07123_ _01370_ _02707_ _02671_ u_arbiter.i_wb_cpu_dbus_sel\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07054_ _02542_ u_cpu.rf_ram.rdata\[4\] _02656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06005_ _01621_ _01622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_82_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07527__I _03004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[53\]_SE net561 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07917__A2 _03254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05928__A1 u_arbiter.i_wb_cpu_dbus_adr\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09119__A1 u_cpu.rf_ram.memory\[36\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07956_ _03291_ _00272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06907_ u_cpu.rf_ram.memory\[136\]\[7\] u_cpu.rf_ram.memory\[137\]\[7\] u_cpu.rf_ram.memory\[138\]\[7\]
+ u_cpu.rf_ram.memory\[139\]\[7\] _01831_ _01832_ _02517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_25_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07887_ u_cpu.rf_ram.memory\[74\]\[2\] _03245_ _03246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08342__A2 _03526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09626_ _04366_ _04367_ _00867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06838_ _02441_ _02443_ _02445_ _02447_ _01807_ _02448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_16_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09557_ _03132_ _04284_ _04318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_110_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06769_ u_cpu.rf_ram.memory\[40\]\[6\] u_cpu.rf_ram.memory\[41\]\[6\] u_cpu.rf_ram.memory\[42\]\[6\]
+ u_cpu.rf_ram.memory\[43\]\[6\] _01736_ _02103_ _02380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_93_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08508_ _03639_ _00476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09488_ u_cpu.rf_ram.memory\[116\]\[4\] _04262_ _04265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10988__A1 u_cpu.rf_ram.memory\[110\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08439_ _03595_ _03590_ _03597_ _00449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06200__S1 _01816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07853__A1 _03195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06900__I0 u_cpu.rf_ram.memory\[72\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09189__I _03915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11450_ _00154_ net334 u_cpu.rf_ram.memory\[48\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10401_ _04198_ u_cpu.rf_ram.memory\[3\]\[6\] _04972_ _04980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10128__I _04809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11381_ _00085_ net176 u_cpu.rf_ram.memory\[80\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10332_ _04937_ _01003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06959__A3 _02565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09358__A1 _04154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10263_ u_cpu.rf_ram.memory\[30\]\[0\] _04895_ _04896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11165__A1 _05456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12002_ _00685_ net415 u_cpu.rf_ram.memory\[38\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10194_ _04854_ _00948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06267__S1 _01699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10912__A1 _05280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12326__CLK net525 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08581__A2 _03287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout370 net372 net370 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout381 net382 net381 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_115_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout392 net393 net392 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_43_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08333__A2 _03529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08268__I _03484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12476__CLK net234 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07172__I _02751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11350__CLK net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06895__A2 _02500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08097__A1 u_cpu.rf_ram.memory\[29\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09833__A2 _04456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07844__A1 _03186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11717_ _00421_ net417 u_cpu.rf_ram.memory\[53\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10239__S _04848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08892__I0 _03574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12697_ u_cpu.rf_ram_if.wdata1_r\[1\] net140 u_cpu.rf_ram_if.wdata1_r\[0\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07121__B _02699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11648_ _00352_ net215 u_cpu.rf_ram.memory\[60\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11579_ _00283_ net350 u_cpu.rf_ram.memory\[68\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout215_I net219 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07072__A2 _02654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09349__A1 _04145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11156__A1 _05444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08021__A1 _03262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06251__I _01601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10903__A1 _05268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07810_ _03083_ _03197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_26_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08790_ _02786_ _03814_ _03815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07741_ _03084_ _03143_ _03151_ _00197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11744__D _00001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07672_ _03101_ _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_77_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06335__A1 _01830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09411_ _04140_ _04213_ _04215_ _00804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_4_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06623_ u_cpu.rf_ram.memory\[92\]\[4\] u_cpu.rf_ram.memory\[93\]\[4\] u_cpu.rf_ram.memory\[94\]\[4\]
+ u_cpu.rf_ram.memory\[95\]\[4\] _02142_ _01915_ _02236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06430__S1 _01799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06886__A2 _02486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11843__CLK net432 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09342_ _04158_ _04162_ _04171_ _00779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout30_I net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06554_ _01400_ _02167_ _02168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08088__A1 _03342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07810__I _03083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09273_ u_cpu.rf_ram.memory\[34\]\[7\] _04116_ _04127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07835__A1 _03197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06485_ _01675_ _02099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08224_ _03458_ _00373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11993__CLK net259 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09588__A1 u_arbiter.i_wb_cpu_rdt\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08155_ _03415_ _03407_ _03416_ _00346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07106_ _02694_ _02595_ _02695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08260__A1 _03417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08086_ _03368_ _03373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12349__CLK net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07037_ _02613_ _02640_ _02643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11147__A1 u_cpu.rf_ram.memory\[27\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06161__I _01777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09760__A1 _04467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12499__CLK net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08988_ u_cpu.rf_ram.memory\[126\]\[6\] _03938_ _03943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10370__A2 _04962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07939_ _03262_ _03274_ _03280_ _00266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09512__A1 u_cpu.rf_ram.memory\[33\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08315__A2 _03517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10950_ _05331_ _01227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10122__A2 _02705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09609_ u_arbiter.i_wb_cpu_dbus_dat\[19\] _04352_ _04356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10881_ u_cpu.rf_ram.memory\[69\]\[0\] _05290_ _05291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06421__S1 _01780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12620_ _01299_ net51 u_cpu.rf_ram.memory\[26\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08079__A1 _03367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09815__A2 _04514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12551_ _01230_ net135 u_cpu.rf_ram.memory\[10\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07826__A1 u_cpu.rf_ram.memory\[129\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09140__C _04032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11502_ _00206_ net99 u_cpu.rf_ram.memory\[17\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12482_ _01161_ net40 u_cpu.rf_ram.memory\[105\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11433_ _00137_ net326 u_cpu.rf_ram.memory\[51\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08626__I0 _03564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11364_ _00068_ net112 u_cpu.rf_ram.memory\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08251__A1 _03405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06101__I1 u_cpu.rf_ram.memory\[109\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10315_ _04927_ _00996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_113_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11295_ u_cpu.rf_ram.memory\[23\]\[1\] _05548_ _05550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11138__A1 u_cpu.rf_ram.memory\[27\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06071__I _01687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10246_ u_arbiter.i_wb_cpu_dbus_adr\[30\] _02691_ _04883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08003__A1 _03264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08554__A2 _03227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10177_ u_cpu.rf_ram.memory\[31\]\[6\] _04840_ _04845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10361__A2 _02586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06660__S1 _01585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08306__A2 _03514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10321__I _04908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11310__A1 _04511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06707__I3 u_cpu.rf_ram.memory\[119\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06412__S1 _01915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout165_I net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout332_I net335 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06270_ _01703_ _01885_ _01709_ _01886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06246__I _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08490__A1 _03602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07293__A2 _02833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09985__C _04575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08242__A1 _03419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06479__S1 _02092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09990__A1 _03115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08793__A2 _03817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09960_ _04492_ _04659_ _04427_ _04660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06643__I2 u_cpu.rf_ram.memory\[138\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11129__A1 _05444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11396__CLK net302 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08911_ _03828_ _03883_ _03890_ _00628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09891_ u_cpu.rf_ram.memory\[114\]\[7\] _04587_ _04598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08545__A2 _03659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08842_ u_cpu.rf_ram.memory\[131\]\[1\] _03848_ _03850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout78_I net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08773_ u_cpu.rf_ram.memory\[134\]\[1\] _03803_ _03805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05985_ _01601_ _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07724_ _02790_ _02891_ _03141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06308__A1 _01778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10104__A2 _04739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07356__I0 _02867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11301__A1 _02903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07655_ _03060_ _03090_ _03092_ _00170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06403__S1 _01905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06606_ u_cpu.rf_ram.memory\[104\]\[4\] u_cpu.rf_ram.memory\[105\]\[4\] u_cpu.rf_ram.memory\[106\]\[4\]
+ u_cpu.rf_ram.memory\[107\]\[4\] _02005_ _01892_ _02219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_13_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12021__CLK net481 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07586_ _02994_ _03036_ _03043_ _00150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_90_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09325_ _04160_ _04162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_40_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07808__A1 u_cpu.rf_ram.memory\[119\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06537_ _01632_ _02151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09256_ _04116_ _04117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06156__I _01685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08481__A1 _03593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06468_ u_cpu.rf_ram.memory\[16\]\[3\] u_cpu.rf_ram.memory\[17\]\[3\] u_cpu.rf_ram.memory\[18\]\[3\]
+ u_cpu.rf_ram.memory\[19\]\[3\] _01852_ _01968_ _02082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_103_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08207_ u_cpu.rf_ram.memory\[19\]\[7\] _03438_ _03449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12171__CLK net386 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09187_ u_cpu.rf_ram.memory\[90\]\[5\] _04064_ _04071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06399_ _01648_ _02014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05995__I _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10415__I0 _04194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09467__I _03912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11739__CLK net152 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08138_ u_cpu.rf_ram.memory\[62\]\[7\] _03393_ _03404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08233__A1 _03410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09981__A1 _04420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08784__A2 _03806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08069_ _03345_ _03356_ _03362_ _00314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10406__I _04982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06634__I2 u_cpu.rf_ram.memory\[70\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10100_ _04701_ _04700_ _04785_ _04459_ _04786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__10591__A2 _05104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11080_ _05361_ _05405_ _05412_ _01276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10031_ _04549_ _04561_ _04725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09733__A1 _04416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08536__A2 _03656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06759__C _01784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10141__I _02756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11982_ _00672_ net411 u_cpu.rf_ram.memory\[123\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05770__A2 _01389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10933_ u_cpu.rf_ram.memory\[59\]\[5\] _05318_ _05322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10864_ u_cpu.rf_ram.memory\[108\]\[3\] _05276_ _05279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12603_ _01282_ net374 u_cpu.cpu.genblk3.csr.mcause3_0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10795_ _05204_ _05232_ _05235_ _01168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12514__CLK net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06158__S0 _01773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08472__A1 _03604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06066__I _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12534_ _01213_ net276 u_cpu.rf_ram.memory\[84\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07275__A2 _02822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_scanchain_local.scan_flop\[56\] u_scanchain_local.module_data_in\[55\] net561 u_arbiter.o_wb_cpu_adr\[18\]
+ net30 u_scanchain_local.module_data_in\[56\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__05825__A3 _01464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12465_ _01144_ net44 u_cpu.rf_ram.memory\[99\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09377__I _02863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11416_ _00120_ net225 u_cpu.rf_ram.memory\[45\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12396_ _01075_ net199 u_cpu.rf_ram.memory\[95\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10031__A1 _04549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11347_ _00051_ net69 u_cpu.rf_ram.memory\[18\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06625__I2 u_cpu.rf_ram.memory\[90\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11278_ u_cpu.rf_ram.memory\[89\]\[2\] _05539_ _05540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06881__S1 _01699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09724__A1 _01438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08527__A2 _03647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10229_ u_arbiter.i_wb_cpu_dbus_adr\[23\] u_arbiter.i_wb_cpu_dbus_adr\[22\] _04873_
+ _04874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10334__A2 _04936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05770_ u_cpu.cpu.immdec.imm24_20\[3\] _01389_ _01421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05761__A2 _01411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10098__A1 _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10986__I _02751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout547_I net550 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07440_ _02900_ _02942_ _02947_ _00100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08456__I _03608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06710__A1 _01647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12194__CLK net403 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07371_ _02745_ _02896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10000__B _04694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09110_ _03977_ _04015_ _04020_ _00697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06322_ _01802_ _01937_ _01805_ _01938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_17_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09041_ _03975_ _03972_ _03976_ _00672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06253_ u_cpu.rf_ram.memory\[60\]\[1\] u_cpu.rf_ram.memory\[61\]\[1\] u_cpu.rf_ram.memory\[62\]\[1\]
+ u_cpu.rf_ram.memory\[63\]\[1\] _01639_ _01668_ _01869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_117_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07018__A2 _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08191__I _03438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06184_ _01797_ _01800_ _01801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10022__A1 _02625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06077__I0 u_cpu.rf_ram.memory\[44\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09963__A1 _04528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08766__A2 _03789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06321__S0 _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06777__B2 _02387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09943_ _04601_ _04609_ _04553_ _04645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06872__S1 _01576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09715__A1 _01438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08518__A2 _03644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05764__B u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09874_ _04587_ _04588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07535__I _03006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09191__A2 _04059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08825_ u_cpu.rf_ram.memory\[132\]\[2\] _03839_ _03840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05968_ _01584_ _01585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08756_ u_cpu.rf_ram.memory\[135\]\[2\] _03794_ _03795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05752__A2 _01389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07707_ u_arbiter.i_wb_cpu_dbus_dat\[5\] _03127_ _03128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_2628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05899_ u_arbiter.i_wb_cpu_dbus_adr\[21\] _01481_ _01527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08687_ u_cpu.rf_ram.memory\[137\]\[1\] _03748_ _03751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11411__CLK net224 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07638_ _03078_ _03064_ _03079_ _00166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07569_ u_cpu.rf_ram.memory\[41\]\[7\] _03021_ _03032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09308_ _03906_ _04150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_122_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11561__CLK net258 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08454__A1 _03606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10580_ u_cpu.rf_ram.memory\[28\]\[0\] _05101_ _05102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07257__A2 _02805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12687__CLK net232 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09239_ _04056_ _04105_ _04107_ _00740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12250_ _00933_ net273 u_cpu.rf_ram.memory\[32\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08206__A1 _03421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11201_ _05451_ _05489_ _05494_ _01315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09954__A1 _04419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08757__A2 _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12181_ _00864_ net389 u_arbiter.i_wb_cpu_dbus_dat\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10136__I _02750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06768__A1 _02372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11132_ _05449_ _05446_ _05450_ _01290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_46_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06863__S1 _01768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06083__I3 u_cpu.rf_ram.memory\[39\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09706__A1 _03114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10072__S _01446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11063_ u_cpu.rf_ram.memory\[87\]\[7\] _05391_ _05402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12067__CLK net282 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10014_ _04477_ _04519_ _04709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_48_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09182__A2 _04058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06615__S1 _01905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[1\] u_cpu.cpu.genblk3.csr.i_mtip net552 u_arbiter.o_wb_cpu_we
+ net20 u_arbiter.i_wb_cpu_ack vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__07193__A1 _02741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05743__A2 u_cpu.cpu.state.genblk1.misalign_trap_sync_r vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11965_ _00661_ net465 u_cpu.rf_ram.memory\[125\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10916_ _05284_ _05303_ _05311_ _01213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11904__CLK net458 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11896_ _00592_ net459 u_cpu.rf_ram.memory\[132\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10847_ _05215_ _05258_ _05266_ _01189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_73_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08445__A1 _03600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07248__A2 _02806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10778_ _05206_ _05220_ _05225_ _01161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12517_ _01196_ net203 u_cpu.rf_ram.memory\[108\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08996__A2 _03946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout128_I net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12448_ _01127_ net88 u_cpu.rf_ram.memory\[103\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09945__A1 _04469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10046__I _04737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08748__A2 _03698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12379_ _01058_ net79 u_cpu.rf_ram.memory\[97\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07420__A2 _02929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06854__S1 _02099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout497_I net499 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06940_ u_cpu.cpu.alu.i_rs1 _02549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input2_I io_in[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06871_ _01656_ _02480_ _01587_ _02481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06606__S1 _01892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11434__CLK net327 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05822_ u_arbiter.i_wb_cpu_dbus_adr\[5\] _01461_ _01466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08610_ u_cpu.rf_ram.memory\[143\]\[2\] _03704_ _03705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09590_ u_arbiter.i_wb_cpu_dbus_dat\[13\] _04338_ _04343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06931__A1 u_cpu.cpu.bufreg2.i_cnt_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05753_ _01402_ _01403_ _01404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08541_ u_cpu.rf_ram.memory\[73\]\[2\] _03659_ _03660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08472_ _03604_ _03610_ _03618_ _00461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07487__A2 _02969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07423_ _02913_ _02926_ _02934_ _00096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10491__A1 _05044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07354_ _02864_ u_cpu.rf_ram.memory\[7\]\[4\] _02879_ _02884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07239__A2 _02804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06305_ _01772_ _01920_ _01921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08987__A2 _03935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07285_ u_cpu.rf_ram.memory\[20\]\[0\] _02834_ _02835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06542__S0 _01787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09024_ u_cpu.rf_ram.memory\[124\]\[4\] _03962_ _03965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10794__A2 _05233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06236_ _01621_ _01852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_117_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08739__A2 _03778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06167_ _01427_ _01784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_105_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10546__A2 _05073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07411__A2 _02926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06098_ _01665_ _01715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06845__S1 _01625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09926_ u_cpu.cpu.immdec.imm24_20\[1\] _04630_ _04631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09857_ _04558_ _04559_ _04571_ _04572_ _04573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07175__A1 _02733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08808_ _03503_ _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08911__A2 _03883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09788_ _04509_ _04510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_73_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06773__I1 u_cpu.rf_ram.memory\[37\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08739_ _03755_ _03778_ _03784_ _00562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11750_ _00007_ net254 u_cpu.rf_ram.rdata\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07478__A2 _02969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08675__A1 _03680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10701_ _03165_ _05162_ _05175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11681_ _00385_ net324 u_cpu.rf_ram.memory\[57\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10609__I0 u_arbiter.i_wb_cpu_rdt\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10632_ _04807_ _05130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08824__I _03834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10563_ u_cpu.rf_ram.memory\[96\]\[4\] _05088_ _05091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08978__A2 _03934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06989__A1 _02527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10785__A2 _05224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12302_ _00024_ net496 u_cpu.cpu.ctrl.pc_plus_offset_cy_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06344__I _01787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10494_ u_cpu.rf_ram.memory\[97\]\[2\] _05047_ _05048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09927__A1 u_cpu.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12233_ _00916_ net359 u_cpu.cpu.immdec.imm19_12_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10537__A2 _05072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12164_ _00847_ net390 u_arbiter.i_wb_cpu_dbus_dat\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07402__A2 _02919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06836__S1 _01585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11457__CLK net327 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11115_ _04952_ _02576_ _05438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[19\] u_arbiter.i_wb_cpu_rdt\[16\] net541 u_arbiter.i_wb_cpu_dbus_dat\[13\]
+ net9 u_arbiter.i_wb_cpu_rdt\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_111_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12095_ _00778_ net408 u_cpu.rf_ram.memory\[118\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09155__A2 _04049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11046_ _05391_ _05392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_42_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07705__A3 u_arbiter.i_wb_cpu_dbus_dat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08902__A2 _03882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09390__I _04202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07961__I0 _02864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07124__B _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06519__I _01650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11948_ _00644_ net461 u_cpu.rf_ram.memory\[127\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08666__A1 _03671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10473__A1 _02701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout245_I net246 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11879_ _00575_ net456 u_cpu.rf_ram.memory\[134\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08969__A2 _03923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout412_I net413 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12232__CLK net360 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07070_ _01430_ _02652_ _02666_ _00010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06295__I3 u_cpu.rf_ram.memory\[119\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07641__A2 _03072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06021_ _01571_ _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_126_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11747__D _00004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12382__CLK net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07972_ u_cpu.rf_ram.memory\[68\]\[0\] _03300_ _03301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09711_ _04427_ _04436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_60_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06923_ u_cpu.cpu.branch_op _02532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_25_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09642_ u_arbiter.i_wb_cpu_dbus_dat\[30\] _04378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_68_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout60_I net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06854_ u_cpu.rf_ram.memory\[56\]\[7\] u_cpu.rf_ram.memory\[57\]\[7\] u_cpu.rf_ram.memory\[58\]\[7\]
+ u_cpu.rf_ram.memory\[59\]\[7\] _01729_ _02099_ _02464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06904__A1 _02507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[67\]_CLK net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10700__A2 _05165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06755__I1 u_cpu.rf_ram.memory\[29\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07813__I _03086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05805_ _01451_ _01452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09573_ _04294_ _04331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06785_ _02008_ _02395_ _02396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05736_ _01379_ _01384_ _01385_ _01386_ _01387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_08524_ _03598_ _03643_ _03649_ _00482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08657__A1 _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10464__A1 _02701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08455_ _02966_ _03202_ _03608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07406_ _02921_ _02923_ _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08386_ _03560_ u_cpu.rf_ram.memory\[9\]\[0\] _03562_ _03563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08409__A1 _03285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07337_ u_cpu.rf_ram_if.wdata1_r\[7\] u_cpu.cpu.o_wdata0 _02734_ _02872_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_52_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09676__S _01437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07268_ _02752_ _02818_ _02823_ _00052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09909__A1 _04400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06219_ _01818_ _01824_ _01829_ _01834_ _01835_ _01836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_3_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09007_ _03913_ _03947_ _03954_ _00660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10615__S _05117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07199_ _02741_ _02773_ _02774_ _00032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10519__A2 _05064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11192__A2 _03165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06443__I0 u_cpu.rf_ram.memory\[128\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout530 net534 net530 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout541 net543 net541 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_24_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09909_ _04400_ _04613_ _04614_ _04615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
Xfanout552 net557 net552 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_120_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout563 net564 net563 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_63_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07148__A1 _02701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07699__A2 _02695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08896__A1 _03367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08819__I _03834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12105__CLK net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11802_ _00498_ net369 u_cpu.rf_ram.memory\[71\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08648__A1 u_cpu.rf_ram.memory\[138\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11733_ _00437_ net145 u_cpu.rf_ram.memory\[9\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06783__B _01587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11664_ _00368_ net121 u_cpu.rf_ram.memory\[5\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07871__A2 _03233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10615_ u_arbiter.i_wb_cpu_rdt\[24\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[8\]
+ _05117_ _05121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11595_ _00299_ net251 u_cpu.rf_ram.memory\[66\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06506__S0 _02005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10758__A2 _05207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06074__I _01609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10546_ _05053_ _05073_ _05080_ _01074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10477_ _04545_ _04453_ _05034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12216_ _00899_ net316 u_cpu.rf_ram.memory\[114\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07387__A1 _02907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11183__A2 _05477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12147_ _00830_ net317 u_cpu.rf_ram.memory\[116\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07139__A1 _01658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout195_I net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12078_ _00761_ net319 u_cpu.rf_ram.memory\[117\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11029_ _05347_ _05380_ _05382_ _01255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08729__I _03777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10694__A1 _05142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout362_I net365 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06570_ u_cpu.rf_ram.memory\[4\]\[4\] u_cpu.rf_ram.memory\[5\]\[4\] u_cpu.rf_ram.memory\[6\]\[4\]
+ u_cpu.rf_ram.memory\[7\]\[4\] _01959_ _02071_ _02183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_52_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10446__A1 u_cpu.cpu.immdec.imm11_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09300__A2 _04142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08240_ _03417_ _03461_ _03468_ _00379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_18_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07862__A2 _03230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08171_ _03426_ _03428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10749__A2 _05201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07122_ _01369_ _01372_ _02707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07053_ _02647_ _02654_ _02655_ _00017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_127_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09295__I _03893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06004_ _01620_ _01621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_86_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11772__CLK net514 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05928__A2 _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07955_ _02855_ u_cpu.rf_ram.memory\[6\]\[1\] _03289_ _03291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12128__CLK net405 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06906_ _02496_ _02515_ _01404_ _02516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_46_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07886_ _03240_ _03245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09625_ u_arbiter.i_wb_cpu_rdt\[23\] _04293_ _04359_ u_arbiter.i_wb_cpu_dbus_dat\[23\]
+ _04367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10685__A1 _05130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06837_ _01786_ _02446_ _01795_ _02447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_56_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12278__CLK net532 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09556_ _04289_ _04316_ _04317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09827__B1 _04453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06768_ _02372_ _02374_ _02376_ _02378_ _01427_ _02379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_97_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08507_ _03572_ u_cpu.rf_ram.memory\[13\]\[5\] _03632_ _03639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_70_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05719_ _01369_ _01370_ u_arbiter.i_wb_cpu_dbus_sel\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09487_ _04247_ _04258_ _04264_ _00831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_12_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06699_ _01720_ _02310_ _01663_ _02311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05998__I _01575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08438_ u_cpu.rf_ram.memory\[142\]\[2\] _03596_ _03597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07853__A2 _03217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06900__I1 u_cpu.rf_ram.memory\[73\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08369_ _03491_ _03549_ _03552_ _00424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10400_ _04979_ _01029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11380_ _00084_ net176 u_cpu.rf_ram.memory\[80\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07605__A2 _03052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10331_ u_cpu.cpu.ctrl.o_ibus_adr\[19\] _04936_ _04931_ u_cpu.cpu.ctrl.o_ibus_adr\[20\]
+ _04937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_109_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06959__A4 _02566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09358__A2 _04174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10262_ _04893_ _04895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_12001_ _00684_ net415 u_cpu.rf_ram.memory\[38\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10193_ u_arbiter.i_wb_cpu_dbus_adr\[7\] u_arbiter.i_wb_cpu_dbus_adr\[6\] _04849_
+ _04854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_65_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05919__A2 _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10912__A2 _05302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout360 net362 net360 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_28_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout371 net372 net371 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_8_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06592__A2 _02200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout382 net393 net382 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_47_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout393 net394 net393 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07541__A1 _02994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06069__I _01685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09294__A1 _04074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11645__CLK net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11716_ _00420_ net426 u_cpu.rf_ram.memory\[53\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08284__I _03497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12696_ _01365_ net379 u_cpu.rf_ram_if.rcnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11228__I0 _02872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11647_ _00351_ net215 u_cpu.rf_ram.memory\[60\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11795__CLK net373 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11578_ _00282_ net349 u_cpu.rf_ram.memory\[68\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout110_I net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10529_ u_cpu.rf_ram.memory\[94\]\[7\] _05059_ _05070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout208_I net209 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09349__A2 _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08021__A2 _03324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10903__A2 _05302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07780__A1 u_cpu.rf_ram.memory\[40\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07740_ u_cpu.rf_ram.memory\[16\]\[6\] _03146_ _03151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07363__I _02888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12420__CLK net264 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07671_ _02831_ _02850_ _03101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_38_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07532__A1 _02980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06335__A2 _01950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09410_ u_cpu.rf_ram.memory\[112\]\[0\] _04214_ _04215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06622_ _01647_ _02225_ _02234_ _02235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_52_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06886__A3 _02495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06553_ u_cpu.rf_ram.memory\[136\]\[3\] u_cpu.rf_ram.memory\[137\]\[3\] u_cpu.rf_ram.memory\[138\]\[3\]
+ u_cpu.rf_ram.memory\[139\]\[3\] _01814_ _01942_ _02167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09341_ u_cpu.rf_ram.memory\[118\]\[7\] _04160_ _04171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08088__A2 _03369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout23_I net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09272_ _04072_ _04118_ _04126_ _00754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06484_ _01671_ _02098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07835__A2 _03205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08223_ _02870_ u_cpu.rf_ram.memory\[5\]\[6\] _03450_ _03458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09588__A2 _04334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08154_ u_cpu.rf_ram.memory\[61\]\[3\] _03413_ _03416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07599__A1 _02987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07105_ _02693_ _02597_ _02694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08085_ _03340_ _03369_ _03372_ _00320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08260__A2 _03473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07036_ _02606_ _02623_ _02641_ _02642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__06271__B2 _01886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11147__A2 _05452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09753__I _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11518__CLK net321 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09760__A2 _04480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08987_ _03913_ _03935_ _03942_ _00652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07771__A1 u_cpu.rf_ram.memory\[40\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07938_ u_cpu.rf_ram.memory\[75\]\[3\] _03278_ _03280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07869_ u_cpu.rf_ram.memory\[77\]\[3\] _03233_ _03235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11668__CLK net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07523__A1 _03000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06177__I2 u_cpu.rf_ram.memory\[70\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09608_ _04355_ _00861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_95_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10880_ _05288_ _05290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09539_ u_arbiter.i_wb_cpu_rdt\[1\] _04290_ _04302_ _04303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08079__A2 _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11083__A1 u_cpu.rf_ram.memory\[88\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12550_ _01229_ net143 u_cpu.rf_ram.memory\[10\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07826__A2 _03208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11501_ _00205_ net106 u_cpu.rf_ram.memory\[17\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10830__A1 _04091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12481_ _01160_ net48 u_cpu.rf_ram.memory\[105\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11432_ _00136_ net368 u_cpu.rf_ram.memory\[51\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11363_ _00067_ net114 u_cpu.rf_ram.memory\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08251__A2 _03473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06101__I2 u_cpu.rf_ram.memory\[110\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06262__A1 _01876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10314_ _01495_ _04922_ _04924_ u_cpu.cpu.ctrl.o_ibus_adr\[13\] _04927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_113_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11294_ _02888_ _05547_ _05549_ _01353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11138__A2 _05452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09200__A1 _02549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10245_ u_arbiter.i_wb_cpu_dbus_adr\[31\] _04882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08003__A2 _03312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10346__B1 _04945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12443__CLK net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10176_ _04827_ _04837_ _04844_ _00940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10897__A1 _05286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08279__I _03493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout190 net191 net190 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_43_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06317__A2 _01931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07514__A1 _02994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout158_I net269 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11074__A1 _05354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[43\]_SE net559 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10821__A1 _05209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout325_I net328 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08490__A2 _03622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12679_ _01357_ net96 u_cpu.rf_ram.memory\[23\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06891__I3 u_cpu.rf_ram.memory\[83\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08242__A2 _03462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09990__A2 u_arbiter.i_wb_cpu_rdt\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08910_ u_cpu.rf_ram.memory\[22\]\[5\] _03886_ _03890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09890_ _04253_ _04589_ _04597_ _00901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09573__I _04294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08841_ _03813_ _03847_ _03849_ _00599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07753__A1 _03071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10512__I _05059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08772_ _03745_ _03802_ _03804_ _00575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05984_ _01407_ _01416_ _01601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07723_ _03135_ _03140_ _00190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_113_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11301__A2 _05547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08917__I _03893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07654_ u_cpu.rf_ram.memory\[50\]\[0\] _03091_ _03092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10360__I0 _02612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06865__C _01733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06605_ _02117_ _02217_ _02218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07585_ u_cpu.rf_ram.memory\[43\]\[4\] _03040_ _03043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09324_ _04160_ _04161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11065__A1 _05300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06536_ _01609_ _02150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09255_ _02722_ _02965_ _04116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06467_ _01596_ _02081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08481__A2 _03621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08206_ _03421_ _03440_ _03448_ _00365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09186_ _03912_ _04070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06398_ _02003_ _02007_ _02010_ _02012_ _01900_ _02013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__05834__A4 _01464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08137_ _03351_ _03395_ _03403_ _00341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08233__A2 _03461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10040__A2 _02530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09981__A2 _04492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08068_ u_cpu.rf_ram.memory\[64\]\[3\] _03360_ _03362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06634__I3 u_cpu.rf_ram.memory\[71\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07019_ u_cpu.cpu.immdec.imm31 _02539_ _02625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__10328__B1 _04931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10030_ _04721_ _04722_ _04723_ _04419_ _04724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_27_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09733__A2 _04418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06547__A2 _02160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08099__I _03004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11981_ _00671_ net410 u_cpu.rf_ram.memory\[123\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10932_ _05280_ _05314_ _05321_ _01219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[66\]_SE net554 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10863_ _04820_ _05278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_77_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09859__S _01446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12602_ _01281_ net373 u_cpu.cpu.genblk3.csr.mcause3_0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11056__A1 _05357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10794_ u_cpu.rf_ram.memory\[106\]\[1\] _05233_ _05235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06158__S1 _01774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12533_ _01212_ net276 u_cpu.rf_ram.memory\[84\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08472__A2 _03610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08562__I _03493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12464_ _01143_ net44 u_cpu.rf_ram.memory\[99\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11415_ _00119_ net224 u_cpu.rf_ram.memory\[45\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xu_scanchain_local.scan_flop\[49\] u_scanchain_local.module_data_in\[48\] net558 u_arbiter.o_wb_cpu_adr\[11\]
+ net28 u_scanchain_local.module_data_in\[49\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
X_12395_ _01074_ net198 u_cpu.rf_ram.memory\[95\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09421__A1 u_cpu.rf_ram.memory\[112\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07178__I _02756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06235__A1 _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10031__A2 _04561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06082__I _01667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11346_ _00050_ net98 u_cpu.rf_ram.memory\[18\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06625__I3 u_cpu.rf_ram.memory\[91\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11833__CLK net478 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11277_ _05534_ _05539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10228_ _02690_ _04873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_80_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07735__A1 _03075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10159_ u_cpu.rf_ram.memory\[32\]\[7\] _04809_ _04834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11983__CLK net410 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout275_I net281 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10098__A2 _04750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout442_I net449 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06710__A2 _02312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06257__I _01678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07370_ _02889_ _02893_ _02895_ _00082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06321_ u_cpu.rf_ram.memory\[76\]\[1\] u_cpu.rf_ram.memory\[77\]\[1\] u_cpu.rf_ram.memory\[78\]\[1\]
+ u_cpu.rf_ram.memory\[79\]\[1\] _01582_ _01803_ _01937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_108_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08463__A2 _03613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09568__I _04318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11363__CLK net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09040_ u_cpu.rf_ram.memory\[123\]\[1\] _03973_ _03976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06252_ _01656_ _01866_ _01867_ _01868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__12489__CLK net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10270__A2 _04898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06183_ u_cpu.rf_ram.memory\[72\]\[0\] u_cpu.rf_ram.memory\[73\]\[0\] u_cpu.rf_ram.memory\[74\]\[0\]
+ u_cpu.rf_ram.memory\[75\]\[0\] _01798_ _01799_ _01800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_11_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07088__I _02633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09963__A2 _04484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06321__S1 _01803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09942_ _04642_ _04638_ _04643_ _04520_ _04644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_67_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout90_I net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05764__C _01378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09873_ _02722_ _04224_ _04587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08824_ _03834_ _03839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08755_ _03789_ _03794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05967_ _01575_ _01584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09479__A1 u_cpu.rf_ram.memory\[116\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07706_ u_arbiter.i_wb_cpu_dbus_dat\[4\] _03126_ _03127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08686_ _03490_ _03750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05898_ u_cpu.cpu.ctrl.o_ibus_adr\[21\] _01525_ _01526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07637_ u_cpu.rf_ram.memory\[47\]\[4\] _03072_ _03079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11038__A1 _05359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06167__I _01427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07568_ _02998_ _03023_ _03031_ _00144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09307_ _04147_ _04142_ _04149_ _00766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06519_ _01650_ _02133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_139_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08454__A2 _03591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07499_ _02983_ _02985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09238_ u_cpu.rf_ram.memory\[35\]\[0\] _04106_ _04107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09169_ _04057_ _04058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08206__A2 _03440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11200_ u_cpu.rf_ram.memory\[24\]\[2\] _05493_ _05494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06217__A1 _01830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10013__A2 _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12180_ _00863_ net388 u_arbiter.i_wb_cpu_dbus_dat\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09954__A2 _04514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06768__A2 _02374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11131_ u_cpu.rf_ram.memory\[27\]\[1\] _05447_ _05450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09706__A2 u_arbiter.i_wb_cpu_rdt\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11062_ _05363_ _05393_ _05401_ _01269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10013_ _04504_ _04701_ _04538_ _04707_ _04503_ _04708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_118_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07193__A2 _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05743__A3 _01393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11964_ _00660_ net465 u_cpu.rf_ram.memory\[125\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10915_ u_cpu.rf_ram.memory\[84\]\[6\] _05306_ _05311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09890__A1 _04253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11895_ _00591_ net456 u_cpu.rf_ram.memory\[132\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11029__A1 _05347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11386__CLK net220 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10846_ u_cpu.rf_ram.memory\[83\]\[6\] _05261_ _05266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08445__A2 _03590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10777_ u_cpu.rf_ram.memory\[105\]\[2\] _05224_ _05225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06456__A1 _01580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12516_ _01195_ net197 u_cpu.rf_ram.memory\[108\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06000__S0 _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08292__I _03503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10252__A2 u_cpu.cpu.state.o_cnt_r\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12447_ _01126_ net77 u_cpu.rf_ram.memory\[102\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11201__A1 _05451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12378_ _01057_ net79 u_cpu.rf_ram.memory\[97\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11329_ _00033_ net217 u_cpu.rf_ram.memory\[82\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12011__CLK net425 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07636__I _03077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout392_I net393 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06870_ u_cpu.rf_ram.memory\[104\]\[7\] u_cpu.rf_ram.memory\[105\]\[7\] u_cpu.rf_ram.memory\[106\]\[7\]
+ u_cpu.rf_ram.memory\[107\]\[7\] _01657_ _01660_ _02480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_39_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05821_ _01463_ _01464_ _01465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12161__CLK net497 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06931__A2 u_cpu.cpu.immdec.imm31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08540_ _03654_ _03659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05752_ u_cpu.cpu.immdec.imm24_20\[4\] _01389_ _01403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07371__I _02745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08133__A1 _03347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08471_ u_cpu.rf_ram.memory\[141\]\[6\] _03613_ _03618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08684__A2 _03748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09881__A1 u_cpu.rf_ram.memory\[114\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07422_ u_cpu.rf_ram.memory\[78\]\[6\] _02929_ _02934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07353_ _02883_ _00077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09298__I _04141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06304_ u_cpu.rf_ram.memory\[80\]\[1\] u_cpu.rf_ram.memory\[81\]\[1\] u_cpu.rf_ram.memory\[82\]\[1\]
+ u_cpu.rf_ram.memory\[83\]\[1\] _01773_ _01774_ _01920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_137_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07284_ _02832_ _02834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_40_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06542__S1 _02040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09023_ _03907_ _03958_ _03964_ _00666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06235_ _01611_ _01850_ _01851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06166_ _01778_ _01781_ _01782_ _01783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07947__A1 _03270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06097_ _01566_ _01608_ _01646_ _01713_ _01714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_28_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09925_ _04481_ _04630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12504__CLK net185 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09856_ _04397_ _04572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08372__A1 _03494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07175__A2 _02752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08807_ _03826_ _03816_ _03827_ _00587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09787_ _04442_ _04509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_2_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06999_ _02584_ _02604_ _02605_ _02593_ _02606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_3138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11259__A1 _02899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08738_ u_cpu.rf_ram.memory\[136\]\[3\] _03782_ _03784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08124__A1 _03335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07281__I _02830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12654__CLK net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08669_ _03673_ _03734_ _03739_ _00537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09872__A1 _02562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10700_ _05148_ _05165_ _05174_ _01134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06230__S0 _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11680_ _00384_ net313 u_cpu.rf_ram.memory\[57\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10609__I1 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10631_ _05129_ _01110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09624__A1 u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06438__A1 _02025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10562_ _05049_ _05084_ _05090_ _01080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_127_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12301_ _00983_ net90 u_cpu.rf_ram.memory\[30\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10493_ _05040_ _05047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_120_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12034__CLK net319 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12232_ _00915_ net360 u_cpu.cpu.immdec.imm7 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12163_ _00846_ net498 u_arbiter.i_wb_cpu_dbus_dat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11114_ _05434_ _05436_ _05437_ _01285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_81_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12094_ _00777_ net408 u_cpu.rf_ram.memory\[118\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12184__CLK net389 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11045_ _05300_ _02877_ _05391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09671__I _04395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07166__A2 _02741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08363__A1 _02831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07705__A4 u_arbiter.i_wb_cpu_dbus_dat\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.output_buffers\[3\]_I net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10170__A1 _04817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06764__I2 u_cpu.rf_ram.memory\[62\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08287__I _02761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07191__I _02767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08115__A1 _03349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11947_ _00643_ net444 u_cpu.rf_ram.memory\[127\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09863__A1 _04458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08666__A2 _03734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06677__A1 _01725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10473__A2 _05004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11878_ _00574_ net510 u_cpu.rf_ram.memory\[135\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout140_I net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10829_ _05217_ _05246_ _05255_ _01182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout238_I net240 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09091__A2 _04007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout405_I net406 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06020_ _01596_ _01637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08750__I _03789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11401__CLK net294 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12527__CLK net339 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06452__I1 u_cpu.rf_ram.memory\[9\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07971_ _03298_ _03300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06601__B2 _02213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10006__B _04615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09710_ _04416_ _04419_ _04434_ _04435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_60_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06922_ _01410_ _02531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_68_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11551__CLK net250 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08354__A1 _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12677__CLK net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09641_ _04376_ _04371_ _04377_ _00872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06853_ _01725_ _02462_ _02463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10161__A1 _03367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05804_ _01450_ _01451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09572_ u_arbiter.i_wb_cpu_dbus_dat\[8\] _04329_ _04330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout53_I net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06784_ u_cpu.rf_ram.memory\[100\]\[6\] u_cpu.rf_ram.memory\[101\]\[6\] u_cpu.rf_ram.memory\[102\]\[6\]
+ u_cpu.rf_ram.memory\[103\]\[6\] _02122_ _01576_ _02395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08106__A1 _03340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08523_ u_cpu.rf_ram.memory\[72\]\[3\] _03647_ _03649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05735_ u_cpu.cpu.state.genblk1.misalign_trap_sync_r _01386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_110_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09854__A1 _04486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09854__B2 _04468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06668__A1 _01590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10464__A2 _04630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08454_ _03606_ _03591_ _03607_ _00454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07405_ _02922_ _02923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_17_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08385_ _03561_ _03562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08409__A2 _03062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05891__A2 _01512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07336_ _02871_ _00072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06445__I _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06515__S1 _01737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07093__A1 _02549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07267_ u_cpu.rf_ram.memory\[18\]\[2\] _02822_ _02823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09006_ u_cpu.rf_ram.memory\[125\]\[5\] _03950_ _03954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06840__A1 _02078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06218_ _01405_ _01835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_121_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07198_ u_cpu.rf_ram.memory\[82\]\[6\] _02753_ _02774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06149_ _01671_ _01766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08593__A1 u_cpu.rf_ram.memory\[70\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06180__I _01683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06443__I1 u_cpu.rf_ram.memory\[129\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout520 net521 net520 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_28_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout531 net534 net531 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_99_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout542 net546 net542 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09908_ _04399_ _04527_ _04614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout553 net557 net553 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout564 net565 net564 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_101_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09393__I0 _04188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09839_ _04544_ _04551_ _04554_ _04555_ _04556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_8_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10152__A1 _04827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08896__A2 _03287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10430__I _04992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11801_ _00497_ net368 u_cpu.rf_ram.memory\[71\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08648__A2 _03726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06659__A1 _01958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11732_ _00436_ net135 u_cpu.rf_ram.memory\[9\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11663_ _00367_ net111 u_cpu.rf_ram.memory\[5\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10614_ _05120_ _01102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06355__I _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11594_ _00298_ net246 u_cpu.rf_ram.memory\[66\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09073__A2 _03995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06506__S1 _01892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10545_ u_cpu.rf_ram.memory\[95\]\[5\] _05076_ _05080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08820__A2 _03836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06831__A1 _01637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10476_ _05033_ _01051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xu_scanchain_local.scan_flop\[31\] u_arbiter.i_wb_cpu_rdt\[28\] net547 u_arbiter.i_wb_cpu_dbus_dat\[25\]
+ net17 u_arbiter.i_wb_cpu_rdt\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
X_12215_ _00898_ net316 u_cpu.rf_ram.memory\[114\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08584__A1 u_cpu.rf_ram.memory\[70\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07387__A2 _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11574__CLK net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06090__I _01706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12146_ _00829_ net397 u_cpu.rf_ram.memory\[116\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12077_ _00760_ net310 u_cpu.rf_ram.memory\[117\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08336__A1 _03501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11028_ u_cpu.rf_ram.memory\[111\]\[0\] _05381_ _05382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10143__A1 u_cpu.rf_ram.memory\[32\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout188_I net191 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05945__I0 u_arbiter.i_wb_cpu_dbus_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout355_I net356 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10446__A2 _04636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout522_I net536 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08170_ _03426_ _03427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07121_ _01394_ _02706_ _02699_ u_cpu.cpu.o_wen0 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_31_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07052_ _02650_ u_cpu.rf_ram_if.rdata1\[3\] _02655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_12_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06822__A1 _01830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11917__CLK net458 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06003_ _01571_ _01620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07378__A2 _02901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10382__A1 _04827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07954_ _03290_ _00271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06681__S0 _01736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08327__A1 _03485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09375__I0 _04192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06905_ _01565_ _02505_ _02514_ _02515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_25_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07885_ _03186_ _03241_ _03244_ _00248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10134__A1 u_cpu.rf_ram.memory\[32\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08878__A2 _02982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09624_ u_arbiter.i_wb_cpu_dbus_dat\[24\] _04319_ _04366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06836_ u_cpu.rf_ram.memory\[0\]\[7\] u_cpu.rf_ram.memory\[1\]\[7\] u_cpu.rf_ram.memory\[2\]\[7\]
+ u_cpu.rf_ram.memory\[3\]\[7\] _02074_ _01585_ _02446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06433__S0 _02047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09555_ u_arbiter.i_wb_cpu_dbus_dat\[4\] _03126_ _04316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09827__A1 _04412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06767_ _02098_ _02377_ _01695_ _02378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09827__B2 _04427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06884__B _01709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08506_ _03638_ _00475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05718_ u_cpu.cpu.bufreg.lsb\[1\] _01370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_19_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09486_ u_cpu.rf_ram.memory\[116\]\[3\] _04262_ _04264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06698_ u_cpu.rf_ram.memory\[96\]\[5\] u_cpu.rf_ram.memory\[97\]\[5\] u_cpu.rf_ram.memory\[98\]\[5\]
+ u_cpu.rf_ram.memory\[99\]\[5\] _02125_ _01693_ _02310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_51_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08437_ _03589_ _03596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_11_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11447__CLK net300 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05864__A2 _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06175__I _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08368_ u_cpu.rf_ram.memory\[52\]\[1\] _03550_ _03552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07319_ _02858_ u_cpu.rf_ram.memory\[1\]\[2\] _02852_ _02859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08299_ _02776_ _03509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11597__CLK net251 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10330_ _04905_ _04936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06813__A1 _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10425__I _04992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10261_ _04893_ _04894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_106_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12000_ _00683_ net401 u_cpu.rf_ram.memory\[38\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07369__A2 _02894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10192_ _04853_ _00947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10373__A1 _04814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06672__S0 _01863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout350 net354 net350 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__08318__A1 _03504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout361 net362 net361 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__09366__I0 _04184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout372 net375 net372 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout383 net384 net383 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_86_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout394 net395 net394 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_19_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08869__A2 _03863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07541__A2 _03007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09818__A1 _04493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11715_ _00419_ net427 u_cpu.rf_ram.memory\[53\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12695_ u_cpu.rf_ram_if.rtrig0 net260 u_cpu.rf_ram_if.rtrig1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12372__CLK net343 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06085__I _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11646_ _00350_ net189 u_cpu.rf_ram.memory\[61\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11577_ _00281_ net347 u_cpu.rf_ram.memory\[68\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07909__I _03253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06804__A1 _02147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[66\]_CLK net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10528_ _05055_ _05061_ _05069_ _01067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout103_I net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10459_ _04692_ _04433_ _04491_ _04514_ _05017_ _05018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_83_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08557__A1 u_cpu.rf_ram.memory\[71\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12129_ _00812_ net410 u_cpu.rf_ram.memory\[122\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06663__S0 _01849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08309__A1 _03491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07644__I _03083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07780__A2 _03172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout472_I net473 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06415__S0 _02029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07670_ _03087_ _03091_ _03100_ _00177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_93_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07532__A2 _03007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06621_ _02227_ _02229_ _02231_ _02233_ _02139_ _02234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_37_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09809__A1 _04526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09340_ _04156_ _04162_ _04170_ _00778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06552_ _02141_ _02165_ _01810_ _02166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[19\]_CLK net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09271_ u_cpu.rf_ram.memory\[34\]\[6\] _04121_ _04126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07296__A1 u_cpu.rf_ram.memory\[20\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06483_ _01666_ _02096_ _02097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08222_ _03457_ _00372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout16_I net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09037__A2 _03973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08153_ _03074_ _03415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07104_ u_cpu.cpu.genblk3.csr.o_new_irq _02693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07599__A2 _03048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08084_ u_cpu.rf_ram.memory\[29\]\[1\] _03370_ _03372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10245__I u_arbiter.i_wb_cpu_dbus_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07035_ _02613_ _02624_ _02640_ _02641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_103_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08548__A1 _03602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07220__A1 u_cpu.rf_ram.memory\[21\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06654__S0 _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08986_ u_cpu.rf_ram.memory\[126\]\[5\] _03938_ _03942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07937_ _03259_ _03274_ _03279_ _00265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10107__A1 _04550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10658__A2 _05131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07868_ _03188_ _03229_ _03234_ _00241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08720__A1 u_cpu.rf_ram.memory\[49\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07523__A2 _02985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06177__I3 u_cpu.rf_ram.memory\[71\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09607_ u_arbiter.i_wb_cpu_rdt\[17\] _04326_ _04321_ u_arbiter.i_wb_cpu_dbus_dat\[17\]
+ _04327_ u_arbiter.i_wb_cpu_dbus_dat\[18\] _04355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_99_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06819_ u_cpu.rf_ram.memory\[136\]\[6\] u_cpu.rf_ram.memory\[137\]\[6\] u_cpu.rf_ram.memory\[138\]\[6\]
+ u_cpu.rf_ram.memory\[139\]\[6\] _01831_ _01832_ _02430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_3_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07799_ u_cpu.rf_ram.memory\[119\]\[2\] _03189_ _03190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09538_ _04297_ _04299_ _04300_ _04301_ _04302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_71_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08385__I _03561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07287__A1 u_cpu.rf_ram.memory\[20\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09469_ _04251_ _04240_ _04252_ _00825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_125_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11500_ _00204_ net106 u_cpu.rf_ram.memory\[17\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12480_ _01159_ net48 u_cpu.rf_ram.memory\[105\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10830__A2 _03310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09028__A2 _03962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11431_ _00135_ net368 u_cpu.rf_ram.memory\[51\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08787__A1 _03763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11362_ _00066_ net112 u_cpu.rf_ram.memory\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10594__A1 _05055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10313_ _04926_ _00995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_98_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06262__A2 _01877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06893__S0 _01752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11293_ u_cpu.rf_ram.memory\[23\]\[0\] _05548_ _05549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_u_scanchain_local.scan_flop\[4\]_D u_arbiter.i_wb_cpu_rdt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08539__A1 _03593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10244_ _04881_ _00971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10346__A1 u_cpu.cpu.ctrl.o_ibus_adr\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06645__S0 _02169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10175_ u_cpu.rf_ram.memory\[31\]\[5\] _04840_ _04844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10897__A2 _05290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout180 net183 net180 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__11612__CLK net238 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout191 net192 net191 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__10649__A2 _05138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07514__A2 _02984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08711__A1 u_cpu.rf_ram.memory\[49\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08295__I _02771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11762__CLK net490 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07278__A1 _02778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10821__A2 _05245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12678_ _01356_ net95 u_cpu.rf_ram.memory\[23\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12118__CLK net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout220_I net221 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11629_ _00333_ net181 u_cpu.rf_ram.memory\[63\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05868__B _01455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout318_I net322 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07639__I _02767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10585__A1 u_cpu.rf_ram.memory\[28\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07450__A1 _02916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12268__CLK net521 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06699__B _01663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08840_ u_cpu.rf_ram.memory\[131\]\[0\] _03848_ _03849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06636__S0 _01934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10888__A2 _05293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07753__A2 _03154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08771_ u_cpu.rf_ram.memory\[134\]\[0\] _03803_ _03804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05764__A1 _01413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05983_ u_cpu.rf_ram.memory\[0\]\[0\] u_cpu.rf_ram.memory\[1\]\[0\] u_cpu.rf_ram.memory\[2\]\[0\]
+ u_cpu.rf_ram.memory\[3\]\[0\] _01598_ _01599_ _01600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07722_ _01821_ _03137_ _03140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_66_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07653_ _03089_ _03091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_65_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10360__I1 _02640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06604_ u_cpu.rf_ram.memory\[108\]\[4\] u_cpu.rf_ram.memory\[109\]\[4\] u_cpu.rf_ram.memory\[110\]\[4\]
+ u_cpu.rf_ram.memory\[111\]\[4\] _02001_ _01717_ _02217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_25_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07584_ _02992_ _03036_ _03042_ _00149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09323_ _03180_ _03286_ _04160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06535_ _02147_ _02148_ _02149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07269__A1 u_cpu.rf_ram.memory\[18\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11065__A2 _03166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09254_ _04074_ _04106_ _04115_ _00747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08933__I _03906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06466_ _02078_ _02079_ _02080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08205_ u_cpu.rf_ram.memory\[19\]\[6\] _03443_ _03448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09185_ _04068_ _04058_ _04069_ _00723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06397_ _01728_ _02011_ _01731_ _02012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_120_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06619__I1 u_cpu.rf_ram.memory\[117\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08136_ u_cpu.rf_ram.memory\[62\]\[6\] _03398_ _03403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06244__A2 _01858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08067_ _03342_ _03356_ _03361_ _00313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07018_ _01374_ _02614_ _02624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09194__A1 _04074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10703__I _05175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06627__S0 _01651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07284__I _02832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07744__A2 _02804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05755__A1 _01404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08969_ _03916_ _03923_ _03931_ _00645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11980_ _00020_ net254 u_cpu.rf_ram_if.rdata1\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11785__CLK net350 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10931_ u_cpu.rf_ram.memory\[59\]\[4\] _05318_ _05321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10862_ _05275_ _05270_ _05277_ _01193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09249__A2 _04109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12601_ _01280_ net374 u_cpu.cpu.genblk3.csr.mcause3_0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11056__A2 _05392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06307__I0 u_cpu.rf_ram.memory\[84\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10793_ _05199_ _05232_ _05234_ _01167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12532_ _01211_ net275 u_cpu.rf_ram.memory\[84\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10803__A2 _05236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12463_ _01142_ net48 u_cpu.rf_ram.memory\[104\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11414_ _00118_ net226 u_cpu.rf_ram.memory\[45\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12394_ _01073_ net198 u_cpu.rf_ram.memory\[95\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12410__CLK net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10567__A1 u_cpu.rf_ram.memory\[96\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11345_ _00049_ net217 u_cpu.rf_ram.memory\[81\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07983__A2 _03303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11276_ _02896_ _05535_ _05538_ _01346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09185__A1 _04068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10227_ _04872_ _00963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12560__CLK net162 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07735__A2 _03142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10158_ _04832_ _04833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_58_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10089_ _04447_ _04775_ _04776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_94_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09488__A2 _04262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[10\]_SE net544 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12687__D u_cpu.rf_ram_if.wdata0_r\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout170_I net172 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06546__I0 u_cpu.rf_ram.memory\[72\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11295__A2 _05548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout268_I net269 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06710__A3 _02321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout435_I net476 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06320_ _01797_ _01935_ _01936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11508__CLK net303 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09660__A2 _04388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06474__A2 _02087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06251_ _01601_ _01867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07671__A1 _02831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12090__CLK net401 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06182_ _01584_ _01799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07423__A1 _02913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06857__S0 _01736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07974__A2 _03300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09941_ _04505_ _04490_ _04643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_98_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08223__I0 _02870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09872_ _02562_ _04398_ _04586_ _00894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout83_I net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08823_ _03819_ _03835_ _03838_ _00592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10730__A1 _05137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08754_ _03750_ _03790_ _03793_ _00568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05966_ _01582_ _01583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08928__I _03902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07705_ _03125_ net36 u_arbiter.i_wb_cpu_dbus_dat\[2\] u_arbiter.i_wb_cpu_dbus_dat\[3\]
+ _03126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XTAP_2608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06876__C _01606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08685_ _03745_ _03747_ _03749_ _00543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05897_ u_cpu.cpu.ctrl.o_ibus_adr\[20\] _01519_ _01525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07636_ _03077_ _03078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[28\]_D u_arbiter.i_wb_cpu_rdt\[25\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11038__A2 _05380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07567_ u_cpu.rf_ram.memory\[41\]\[6\] _03026_ _03031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10097__I0 u_arbiter.i_wb_cpu_rdt\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09306_ u_cpu.rf_ram.memory\[120\]\[2\] _04148_ _04149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09100__A1 _03988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06518_ _01904_ _02131_ _01744_ _02132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_142_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12433__CLK net160 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07498_ _02983_ _02984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_70_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09237_ _04104_ _04106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06304__I3 u_cpu.rf_ram.memory\[83\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06449_ _02055_ _02057_ _02059_ _02063_ _01835_ _02064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XANTENNA__07662__A1 _03075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09695__S _04417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09168_ _02731_ _02938_ _04057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10549__A1 u_cpu.rf_ram.memory\[95\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08119_ _03353_ _03383_ _03392_ _00334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06217__A2 _01833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06848__S0 _01747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09099_ u_cpu.rf_ram.memory\[37\]\[7\] _04002_ _04013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11130_ _02745_ _05449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_79_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11061_ u_cpu.rf_ram.memory\[87\]\[6\] _05396_ _05401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[33\]_SE net550 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10012_ _04505_ _04411_ _04504_ _04707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08914__A1 u_cpu.rf_ram.memory\[22\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05728__A1 u_cpu.cpu.decode.opcode\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10721__A1 _03002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08838__I _03846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09714__I0 u_arbiter.i_wb_cpu_rdt\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11963_ _00659_ net445 u_cpu.rf_ram.memory\[125\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[19\]_D u_arbiter.i_wb_cpu_rdt\[16\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_10914_ _05282_ _05303_ _05310_ _01212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11894_ _00590_ net458 u_cpu.rf_ram.memory\[133\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11029__A2 _05380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10845_ _05213_ _05258_ _05265_ _01188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05900__A1 _01524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10776_ _05219_ _05224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10788__A1 _05217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[61\] u_scanchain_local.module_data_in\[60\] net555 u_arbiter.o_wb_cpu_adr\[23\]
+ net23 u_scanchain_local.module_data_in\[61\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__06456__A2 _02068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12515_ _01194_ net197 u_cpu.rf_ram.memory\[108\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06000__S1 _01616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10608__I _03116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12446_ _01125_ net77 u_cpu.rf_ram.memory\[102\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12377_ _01056_ net74 u_cpu.rf_ram.memory\[97\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06839__S0 _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11328_ _00032_ net204 u_cpu.rf_ram.memory\[82\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09158__A1 _03980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11259_ _02899_ _05523_ _05528_ _01339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08905__A1 _03821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout385_I net388 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10712__A1 _05140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05820_ u_cpu.cpu.genblk1.align.ctrl_misal u_cpu.cpu.ctrl.o_ibus_adr\[4\] u_cpu.cpu.ctrl.o_ibus_adr\[3\]
+ u_cpu.cpu.ctrl.o_ibus_adr\[2\] _01464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XANTENNA__08381__A2 _03548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07652__I _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05751_ u_cpu.cpu.immdec.imm19_12_20\[8\] _01401_ _01402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout552_I net557 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11268__A2 _05522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11174__I _05476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08133__A2 _03394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08470_ _03602_ _03610_ _03617_ _00460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11330__CLK net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12456__CLK net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07421_ _02910_ _02926_ _02933_ _00095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07892__A1 _03193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06695__A2 _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07352_ _02861_ u_cpu.rf_ram.memory\[7\]\[3\] _02879_ _02883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06303_ _01766_ _01918_ _01770_ _01919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_17_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10518__I _05059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07283_ _02832_ _02833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11480__CLK net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06217__B _01419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09022_ u_cpu.rf_ram.memory\[124\]\[3\] _03962_ _03964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06234_ u_cpu.rf_ram.memory\[20\]\[1\] u_cpu.rf_ram.memory\[21\]\[1\] u_cpu.rf_ram.memory\[22\]\[1\]
+ u_cpu.rf_ram.memory\[23\]\[1\] _01849_ _01616_ _01850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_30_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06165_ _01627_ _01782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[56\]_SE net561 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07947__A2 _03275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06096_ _01647_ _01682_ _01712_ _01713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_46_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09924_ _04628_ _04629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09855_ _04560_ _04562_ _04570_ _04571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08372__A2 _03549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08806_ u_cpu.rf_ram.memory\[133\]\[4\] _03822_ _03827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09786_ _04459_ _04507_ _04508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06998_ _01375_ _02605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06383__B2 _01997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08737_ _03752_ _03778_ _03783_ _00561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11259__A2 _05523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06773__I3 u_cpu.rf_ram.memory\[39\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05949_ _01565_ _01566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08124__A2 _03394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06178__I _01627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08668_ u_cpu.rf_ram.memory\[39\]\[2\] _03738_ _03739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09872__A2 _04398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07883__A1 _03179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06230__S1 _01599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06686__A2 _02297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07619_ _03063_ _03065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08599_ u_cpu.rf_ram.memory\[70\]\[7\] _03686_ _03697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10630_ u_arbiter.i_wb_cpu_rdt\[31\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\]
+ _03116_ _05129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09624__A2 _04319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05810__I _01455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10561_ u_cpu.rf_ram.memory\[96\]\[3\] _05088_ _05090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12300_ _00982_ net79 u_cpu.rf_ram.memory\[30\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11973__CLK net446 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10492_ _04816_ _05046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_12231_ _00914_ net383 u_cpu.cpu.immdec.imm30_25\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07938__A2 _03278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12162_ _00845_ net497 u_arbiter.i_wb_cpu_dbus_dat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12329__CLK net504 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11113_ _02576_ _05436_ _04032_ _05437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12093_ _00776_ net404 u_cpu.rf_ram.memory\[118\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07673__S _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11044_ _05365_ _05381_ _05390_ _01262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_49_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08363__A2 _03425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11353__CLK net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12479__CLK net242 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10170__A2 _04836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08115__A2 _03383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06088__I _01704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11946_ _00642_ net444 u_cpu.rf_ram.memory\[127\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07874__A1 _03195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11877_ _00573_ net516 u_cpu.rf_ram.memory\[135\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10828_ u_cpu.rf_ram.memory\[107\]\[7\] _05244_ _05255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06429__A2 _02043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout133_I net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10759_ _05211_ _05201_ _05212_ _01155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_12_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout300_I net304 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12429_ _01108_ net363 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07647__I _02777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08051__A1 _03349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10933__A1 u_cpu.rf_ram.memory\[59\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12205__D _00888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07970_ _03298_ _03299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06601__A2 _02209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06921_ _02529_ _02530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08354__A2 _03537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09640_ u_arbiter.i_wb_cpu_rdt\[28\] _04326_ _04295_ u_arbiter.i_wb_cpu_dbus_dat\[28\]
+ _04377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_68_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06852_ u_cpu.rf_ram.memory\[60\]\[7\] u_cpu.rf_ram.memory\[61\]\[7\] u_cpu.rf_ram.memory\[62\]\[7\]
+ u_cpu.rf_ram.memory\[63\]\[7\] _02095_ _01633_ _02462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_95_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06365__A1 _01656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10161__A2 _03062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05803_ _01432_ u_cpu.cpu.state.ibus_cyc _01450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09571_ _04327_ _04329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06783_ _02004_ _02393_ _01587_ _02394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_110_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09303__A1 _04145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11846__CLK net421 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08522_ _03595_ _03643_ _03648_ _00481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05734_ u_cpu.cpu.genblk3.csr.o_new_irq _01385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_24_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06117__A1 _01719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout46_I net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08453_ u_cpu.rf_ram.memory\[142\]\[7\] _03589_ _03607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07865__A1 _03186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06668__A2 _02279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07404_ _02729_ _02848_ _02922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08384_ _03285_ _03020_ _03561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_91_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11996__CLK net400 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07335_ _02870_ u_cpu.rf_ram.memory\[1\]\[6\] _02851_ _02871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_17_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07617__A1 _03018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08941__I _03912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08290__A1 _03501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07266_ _02817_ _02822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09005_ _03910_ _03946_ _03953_ _00659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06217_ _01830_ _01833_ _01419_ _01834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08417__I0 _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07197_ _02772_ _02773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08042__A1 _03342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06148_ _01761_ _01764_ _01765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10924__A1 u_cpu.rf_ram.memory\[59\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09790__A1 _04416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08593__A2 _03691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09790__B2 _04423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06079_ _01691_ _01694_ _01695_ _01696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11376__CLK net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout510 net511 net510 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_28_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout521 net522 net521 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_09907_ _04443_ _04546_ _04613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout532 net534 net532 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_28_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12621__CLK net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout543 net546 net543 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_58_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout554 net556 net554 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout565 net4 net565 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_101_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09838_ _03118_ _04438_ _04555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08388__I _02854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06356__A1 _01619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05805__I _01451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10152__A2 _04811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09769_ _04478_ _04491_ _04492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_73_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11800_ _00496_ net348 u_cpu.rf_ram.memory\[71\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11731_ _00435_ net132 u_cpu.rf_ram.memory\[9\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06659__A2 _02270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12001__CLK net415 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11662_ _00366_ net182 u_cpu.rf_ram.memory\[19\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10613_ u_arbiter.i_wb_cpu_rdt\[23\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[7\]
+ _05117_ _05120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10158__I _04832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07608__A1 _02996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11593_ _00297_ net244 u_cpu.rf_ram.memory\[66\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10544_ _05051_ _05072_ _05079_ _01073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08281__A1 u_cpu.rf_ram.memory\[56\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12151__CLK net401 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10475_ _05030_ _05032_ _04466_ _05033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06831__A2 _02440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12214_ _00897_ net316 u_cpu.rf_ram.memory\[114\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11719__CLK net332 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08584__A2 _03688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12145_ _00828_ net397 u_cpu.rf_ram.memory\[116\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_scanchain_local.scan_flop\[24\] u_arbiter.i_wb_cpu_rdt\[21\] net541 u_arbiter.i_wb_cpu_dbus_dat\[18\]
+ net9 u_arbiter.i_wb_cpu_rdt\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_68_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08499__S _03633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12076_ _00759_ net318 u_cpu.rf_ram.memory\[117\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11869__CLK net516 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08336__A2 _03525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09533__A1 u_arbiter.i_wb_cpu_dbus_dat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11027_ _05379_ _05381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_42_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05715__I _01367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12695__D u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07847__A1 _03188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout250_I net255 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11929_ _00625_ net419 u_cpu.rf_ram.memory\[22\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout348_I net349 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout515_I net522 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07120_ u_cpu.cpu.immdec.imm11_7\[4\] _02702_ _02704_ _02705_ _02706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_9_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08272__A1 u_cpu.rf_ram.memory\[56\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07051_ _02648_ u_cpu.rf_ram.rdata\[3\] _02654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06822__A2 _02432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11399__CLK net293 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06002_ _01596_ _01619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12644__CLK net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10017__B _04619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09772__A1 _04484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10382__A2 _04962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07953_ _02846_ u_cpu.rf_ram.memory\[6\]\[0\] _03289_ _03290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06681__S1 _02103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08327__A2 _03525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06904_ _02507_ _02509_ _02511_ _02513_ _01711_ _02514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_56_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07884_ u_cpu.rf_ram.memory\[74\]\[1\] _03242_ _03244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10134__A2 _04811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09623_ _04364_ _04365_ _00866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06835_ _01580_ _02444_ _02445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06433__S1 _01803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09554_ _04310_ _04312_ _04314_ _04315_ _00847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08936__I _02761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06766_ u_cpu.rf_ram.memory\[56\]\[6\] u_cpu.rf_ram.memory\[57\]\[6\] u_cpu.rf_ram.memory\[58\]\[6\]
+ u_cpu.rf_ram.memory\[59\]\[6\] _01729_ _02099_ _02377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_36_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09827__A2 _04434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07840__I _03215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05717_ u_cpu.cpu.bufreg.lsb\[0\] _01369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08505_ _03570_ u_cpu.rf_ram.memory\[13\]\[4\] _03633_ _03638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07838__A1 _03033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08886__I0 _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09485_ _04244_ _04258_ _04263_ _00830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06697_ _02008_ _02308_ _02309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08436_ _03493_ _03595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_36_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06510__A1 _02008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12174__CLK net363 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08638__I0 _03576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08367_ _03485_ _03549_ _03551_ _00423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09767__I _04432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07318_ _02857_ _02858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_109_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07066__A2 _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08298_ _03507_ _03488_ _03508_ _00397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07249_ u_cpu.rf_ram.memory\[81\]\[3\] _02810_ _02812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10260_ _03367_ _02921_ _04893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10191_ u_arbiter.i_wb_cpu_dbus_adr\[6\] u_arbiter.i_wb_cpu_dbus_adr\[5\] _04849_
+ _04853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_121_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06121__S0 _01736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10373__A2 _04961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06672__S1 _01748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout340 net345 net340 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout351 net354 net351 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__09515__A1 _04255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08318__A2 _03514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout362 net365 net362 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_93_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09366__I1 u_cpu.rf_ram.memory\[8\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout373 net374 net373 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_43_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout384 net385 net384 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_101_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout395 net539 net395 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_46_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09818__A2 _04477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07829__A1 _03191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12517__CLK net203 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11272__I _05534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11714_ _00418_ net450 u_cpu.rf_ram.memory\[53\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12694_ _01364_ net379 u_cpu.rf_ram_if.rgnt vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11645_ _00349_ net189 u_cpu.rf_ram.memory\[61\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11541__CLK net249 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11576_ _00280_ net340 u_cpu.rf_ram.memory\[68\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10527_ u_cpu.rf_ram.memory\[94\]\[6\] _05064_ _05069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06804__A2 _02414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07197__I _02772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10458_ _04497_ _04509_ _05017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09754__A1 _04475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06407__I2 u_cpu.rf_ram.memory\[118\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10389_ _04184_ u_cpu.rf_ram.memory\[3\]\[0\] _04973_ _04974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_48_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12128_ _00811_ net405 u_cpu.rf_ram.memory\[112\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06663__S1 _01965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout298_I net305 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09506__A1 u_cpu.rf_ram.memory\[33\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08309__A2 _03513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12059_ _00742_ net307 u_cpu.rf_ram.memory\[35\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10116__A2 _04796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12047__CLK net500 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06415__S1 _01768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout465_I net467 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06620_ _01751_ _02232_ _01755_ _02233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_25_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09809__A2 _04479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06551_ _02026_ _02155_ _02164_ _02165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__12197__CLK net396 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09270_ _04070_ _04118_ _04125_ _00753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06276__I _01659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06482_ u_cpu.rf_ram.memory\[60\]\[3\] u_cpu.rf_ram.memory\[61\]\[3\] u_cpu.rf_ram.memory\[62\]\[3\]
+ u_cpu.rf_ram.memory\[63\]\[3\] _02095_ _01668_ _02096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07296__A2 _02837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08221_ _02867_ u_cpu.rf_ram.memory\[5\]\[5\] _03450_ _03457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08152_ _03412_ _03407_ _03414_ _00345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07103_ _01431_ u_cpu.cpu.ctrl.pc_plus_offset_cy_r _02635_ _02692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_140_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08083_ _03335_ _03369_ _03371_ _00319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08796__A2 _03817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06351__S0 _01849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07034_ _02638_ _02586_ _02639_ _02640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08548__A2 _03656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06654__S1 _01838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08985_ _03910_ _03934_ _03941_ _00651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10261__I _04893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07936_ u_cpu.rf_ram.memory\[75\]\[2\] _03278_ _03279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07867_ u_cpu.rf_ram.memory\[77\]\[2\] _03233_ _03234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11414__CLK net226 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09606_ _04353_ _04354_ _00860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06818_ _02409_ _02428_ _01404_ _02429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07798_ _03182_ _03189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09537_ net36 _04288_ _04301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06749_ _01786_ _02359_ _01795_ _02360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06186__I _01706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08484__A1 _03595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11564__CLK net343 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09468_ u_cpu.rf_ram.memory\[115\]\[5\] _04245_ _04252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08419_ _03570_ u_cpu.rf_ram.memory\[15\]\[4\] _03579_ _03584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_36_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09399_ _04194_ u_cpu.rf_ram.memory\[11\]\[4\] _04203_ _04208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06590__S0 _01871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11430_ _00134_ net370 u_cpu.rf_ram.memory\[51\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08236__A1 _03412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11361_ _00065_ net65 u_cpu.rf_ram.memory\[20\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08787__A2 _03803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06798__A1 _01647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10312_ u_cpu.cpu.ctrl.o_ibus_adr\[11\] _04922_ _04924_ _01495_ _04926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_49_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11292_ _05546_ _05548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06893__S1 _02151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09736__A1 _04412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08539__A2 _03655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10243_ u_arbiter.i_wb_cpu_dbus_adr\[30\] u_arbiter.i_wb_cpu_dbus_adr\[29\] _04848_
+ _04881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07211__A2 _02784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10174_ _04824_ _04836_ _04843_ _00939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06645__S1 _01816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05773__A2 _01367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout170 net172 net170 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_43_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07681__S _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout181 net183 net181 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_87_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout192 net193 net192 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_47_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08711__A2 _03767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08475__A1 _02981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07278__A2 _02819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09401__S _04202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06029__C _01428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12677_ _01355_ net95 u_cpu.rf_ram.memory\[23\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06581__S0 _01622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10409__I0 _04188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08227__A1 _02937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11628_ _00332_ net181 u_cpu.rf_ram.memory\[63\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10034__A1 _04721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09975__A1 _04397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08778__A2 _03806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11559_ _00263_ net257 u_cpu.rf_ram.memory\[75\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10585__A2 _05104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06636__S1 _01763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11437__CLK net324 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06261__I0 u_cpu.rf_ram.memory\[40\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08950__A2 _03895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05982_ _01584_ _01599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08770_ _03801_ _03803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05764__A2 _01414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07721_ _03139_ _00189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07652_ _03089_ _03090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11587__CLK net251 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06603_ _01566_ _02187_ _02196_ _02215_ _02216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_20_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07583_ u_cpu.rf_ram.memory\[43\]\[3\] _03040_ _03042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09322_ _04158_ _04143_ _04159_ _00771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06534_ u_cpu.rf_ram.memory\[80\]\[3\] u_cpu.rf_ram.memory\[81\]\[3\] u_cpu.rf_ram.memory\[82\]\[3\]
+ u_cpu.rf_ram.memory\[83\]\[3\] _01773_ _02033_ _02148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08466__A1 _03598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07269__A2 _02822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10273__A1 _04824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09253_ u_cpu.rf_ram.memory\[35\]\[7\] _04104_ _04115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06465_ u_cpu.rf_ram.memory\[20\]\[3\] u_cpu.rf_ram.memory\[21\]\[3\] u_cpu.rf_ram.memory\[22\]\[3\]
+ u_cpu.rf_ram.memory\[23\]\[3\] _01849_ _01965_ _02079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_107_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06572__S0 _02074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08204_ _03419_ _03440_ _03447_ _00364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09184_ u_cpu.rf_ram.memory\[90\]\[4\] _04064_ _04069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06396_ u_cpu.rf_ram.memory\[96\]\[2\] u_cpu.rf_ram.memory\[97\]\[2\] u_cpu.rf_ram.memory\[98\]\[2\]
+ u_cpu.rf_ram.memory\[99\]\[2\] _01729_ _01641_ _02011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_33_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10025__A1 _04713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09966__A1 _02529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08135_ _03349_ _03395_ _03402_ _00340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06619__I2 u_cpu.rf_ram.memory\[118\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08066_ u_cpu.rf_ram.memory\[64\]\[2\] _03360_ _03361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12212__CLK net318 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07441__A2 _02946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09718__A1 _04439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07017_ _02612_ _02615_ _02575_ _02622_ _02623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_89_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10328__A2 _04929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09194__A2 _04059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06627__S1 _02033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[50\]_CLK net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12362__CLK net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08968_ u_cpu.rf_ram.memory\[127\]\[6\] _03926_ _03931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06952__A1 _02559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05755__A2 _01405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07919_ u_cpu.rf_ram.memory\[76\]\[5\] _03260_ _03267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08899_ u_cpu.rf_ram.memory\[22\]\[0\] _03883_ _03884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10930_ _05278_ _05314_ _05320_ _01218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[65\]_CLK net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10500__A2 _05047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10861_ u_cpu.rf_ram.memory\[108\]\[2\] _05276_ _05277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12600_ _01279_ net378 u_cpu.cpu.genblk3.csr.mcause3_0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10792_ u_cpu.rf_ram.memory\[106\]\[0\] _05233_ _05234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10264__A1 _04808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12531_ _01210_ net271 u_cpu.rf_ram.memory\[84\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08209__A1 _02786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12462_ _01141_ net43 u_cpu.rf_ram.memory\[104\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10016__A1 _04680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09957__A1 _04651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11413_ _00117_ net227 u_cpu.rf_ram.memory\[45\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12393_ _01072_ net198 u_cpu.rf_ram.memory\[95\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06315__S0 _01792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10567__A2 _05088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11344_ _00048_ net207 u_cpu.rf_ram.memory\[81\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09709__A1 _04429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06640__B1 _02250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12705__CLK net353 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11275_ u_cpu.rf_ram.memory\[89\]\[1\] _05536_ _05538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10319__A2 _04929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09185__A2 _04058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10226_ u_arbiter.i_wb_cpu_dbus_adr\[22\] u_arbiter.i_wb_cpu_dbus_adr\[21\] _04867_
+ _04872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_u_scanchain_local.scan_flop\[18\]_CLK net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10157_ _02776_ _04832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06943__A1 _02530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10088_ _04401_ _04642_ _04443_ _04774_ _04553_ _04775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_23_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05723__I u_cpu.cpu.decode.opcode\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06546__I1 u_cpu.rf_ram.memory\[73\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout163_I net164 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08448__A1 _03602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout330_I net332 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07120__A1 u_cpu.cpu.immdec.imm11_7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout428_I net429 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06250_ u_cpu.rf_ram.memory\[48\]\[1\] u_cpu.rf_ram.memory\[49\]\[1\] u_cpu.rf_ram.memory\[50\]\[1\]
+ u_cpu.rf_ram.memory\[51\]\[1\] _01657_ _01660_ _01866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__12235__CLK net263 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07671__A2 _02850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10007__A1 _04700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09948__A1 _04629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06181_ _01612_ _01798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_15_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08620__A1 u_cpu.rf_ram.memory\[143\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07423__A2 _02926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06077__I3 u_cpu.rf_ram.memory\[47\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06857__S1 _02103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09940_ _04489_ _04642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07385__I _02906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09871_ _04558_ _04574_ _04584_ _04585_ _04586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07187__A1 _02733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06234__I0 u_cpu.rf_ram.memory\[20\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08822_ u_cpu.rf_ram.memory\[132\]\[1\] _03836_ _03838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08753_ u_cpu.rf_ram.memory\[135\]\[1\] _03791_ _03793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05965_ _01581_ _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07704_ u_arbiter.i_wb_cpu_dbus_dat\[0\] _03125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05896_ _01455_ _01524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08684_ u_cpu.rf_ram.memory\[137\]\[0\] _03748_ _03749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07635_ _02762_ _03077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06793__S0 _02133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08439__A1 _03595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08944__I _02771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07566_ _02996_ _03023_ _03030_ _00143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10246__A1 u_arbiter.i_wb_cpu_dbus_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09305_ _04141_ _04148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09100__A2 _04004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10097__I1 u_arbiter.i_wb_cpu_rdt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06517_ u_cpu.rf_ram.memory\[120\]\[3\] u_cpu.rf_ram.memory\[121\]\[3\] u_cpu.rf_ram.memory\[122\]\[3\]
+ u_cpu.rf_ram.memory\[123\]\[3\] _01741_ _01905_ _02131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_126_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10187__S _04849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07497_ _02965_ _02982_ _02983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10797__A2 _05236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09236_ _04104_ _04105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06464__I _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08880__S _03872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07662__A2 _03090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06448_ _02060_ _02062_ _01419_ _02063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11602__CLK net243 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09167_ _03893_ _04056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06379_ _01706_ _01994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10549__A2 _05071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08118_ u_cpu.rf_ram.memory\[63\]\[7\] _03381_ _03392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08611__A1 _03673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07414__A2 _02929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09098_ _03986_ _04004_ _04012_ _00693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06848__S1 _01748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08049_ _03080_ _03349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11752__CLK net479 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11060_ _05361_ _05393_ _05400_ _01268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10011_ u_arbiter.i_wb_cpu_rdt\[30\] u_arbiter.i_wb_cpu_rdt\[14\] _01447_ _04706_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_103_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08914__A2 _03881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05728__A2 u_cpu.cpu.branch_op vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06925__A1 u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10721__A2 _05162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11962_ _00658_ net445 u_cpu.rf_ram.memory\[125\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08678__A1 u_cpu.rf_ram.memory\[39\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10913_ u_cpu.rf_ram.memory\[84\]\[5\] _05306_ _05310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11893_ _00589_ net468 u_cpu.rf_ram.memory\[133\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06784__S0 _02122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12258__CLK net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10844_ u_cpu.rf_ram.memory\[83\]\[5\] _05261_ _05265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10775_ _05204_ _05220_ _05223_ _01160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_125_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10788__A2 _05221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12514_ _01193_ net196 u_cpu.rf_ram.memory\[108\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08850__A1 _03826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[54\] u_scanchain_local.module_data_in\[53\] net561 u_arbiter.o_wb_cpu_adr\[16\]
+ net29 u_scanchain_local.module_data_in\[54\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
X_12445_ _01124_ net76 u_cpu.rf_ram.memory\[102\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08602__A1 _03061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12376_ _01055_ net79 u_cpu.rf_ram.memory\[97\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06839__S1 _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11327_ _00031_ net170 u_cpu.rf_ram.memory\[82\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05718__I u_cpu.cpu.bufreg.lsb\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10960__A2 _05337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11258_ u_cpu.rf_ram.memory\[100\]\[2\] _05527_ _05528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07169__A1 _02748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10209_ u_arbiter.i_wb_cpu_dbus_adr\[14\] u_arbiter.i_wb_cpu_dbus_adr\[13\] _04861_
+ _04863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08905__A2 _03882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11189_ _05460_ _05478_ _05486_ _01311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10712__A2 _05176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12698__D u_cpu.rf_ram_if.wdata1_r\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout280_I net281 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout378_I net380 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06392__A2 _02006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05750_ _01367_ _01401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08669__A1 _03673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout545_I net546 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07341__A1 _02719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06775__S0 _01767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07420_ u_cpu.rf_ram.memory\[78\]\[5\] _02929_ _02933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07892__A2 _03241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07351_ _02882_ _00076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09094__A1 _03982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11625__CLK net176 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10779__A2 _05224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06302_ u_cpu.rf_ram.memory\[88\]\[1\] u_cpu.rf_ram.memory\[89\]\[1\] u_cpu.rf_ram.memory\[90\]\[1\]
+ u_cpu.rf_ram.memory\[91\]\[1\] _01767_ _01768_ _01918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_52_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06284__I _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07282_ _02790_ _02831_ _02832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08841__A1 _03813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09021_ _03903_ _03958_ _03963_ _00665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06233_ _01573_ _01849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_121_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09809__B _04528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09595__I _04311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11775__CLK net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06164_ u_cpu.rf_ram.memory\[84\]\[0\] u_cpu.rf_ram.memory\[85\]\[0\] u_cpu.rf_ram.memory\[86\]\[0\]
+ u_cpu.rf_ram.memory\[87\]\[0\] _01779_ _01780_ _01781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_121_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06095_ _01690_ _01696_ _01701_ _01710_ _01711_ _01712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_116_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09923_ _04465_ _04627_ _04628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_132_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09854_ _04486_ _04564_ _04569_ _04468_ _04570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07955__I0 _02855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08805_ _03500_ _03826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09785_ _04503_ _04506_ _04457_ _04492_ _04507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_3107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06997_ _02559_ _02587_ _02590_ _02603_ _02604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__06383__A2 _01990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08736_ u_cpu.rf_ram.memory\[136\]\[2\] _03782_ _03783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05948_ _01420_ _01421_ _01565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09857__B1 _04571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10467__A1 _04692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09321__A2 _04141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08667_ _03733_ _03738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05879_ _01451_ _01512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_14_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06766__S0 _01729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07618_ _03063_ _03064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07883__A2 _03241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08598_ _03682_ _03688_ _03696_ _00509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07549_ _02782_ _02936_ _03019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__09085__A1 _03969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10560_ _05046_ _05084_ _05089_ _01079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08832__A1 _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09219_ _04056_ _04093_ _04095_ _00732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10491_ _05044_ _05041_ _05045_ _01054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12230_ _00913_ net361 u_cpu.cpu.immdec.imm30_25\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07399__A1 _02916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12161_ _00844_ net497 u_arbiter.i_wb_cpu_dbus_dat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11112_ _02566_ _04030_ _05435_ _05436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_1_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12092_ _00775_ net404 u_cpu.rf_ram.memory\[118\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11043_ u_cpu.rf_ram.memory\[111\]\[7\] _05379_ _05390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08899__A1 u_cpu.rf_ram.memory\[22\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06797__C _02139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10458__A1 _04497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11945_ _00641_ net444 u_cpu.rf_ram.memory\[127\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06757__S0 _01622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07874__A2 _03230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11876_ _00572_ net516 u_cpu.rf_ram.memory\[135\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10619__I _03116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10827_ _05215_ _05246_ _05254_ _01181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09076__A1 _03984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06509__S0 _02122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11798__CLK net368 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10758_ u_cpu.rf_ram.memory\[79\]\[4\] _05207_ _05212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08823__A1 _03819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06685__I0 u_cpu.rf_ram.memory\[36\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout126_I net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10689_ u_cpu.rf_ram.memory\[103\]\[2\] _05168_ _05169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12428_ _01107_ net364 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11186__A2 _05481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08051__A2 _03338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12359_ _01038_ net138 u_cpu.rf_ram.memory\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10933__A2 _05318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout495_I net499 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06988__B _01374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06920_ _02528_ _02529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09000__A1 u_cpu.rf_ram.memory\[125\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12423__CLK net357 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07011__B1 u_cpu.cpu.mem_bytecnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06851_ _01569_ _02460_ _01602_ _02461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_68_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07562__A1 _02992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06365__A2 _01979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06500__C _01711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05802_ _01434_ _01448_ _01449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09570_ _04328_ _00850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_95_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06279__I _01667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06782_ u_cpu.rf_ram.memory\[104\]\[6\] u_cpu.rf_ram.memory\[105\]\[6\] u_cpu.rf_ram.memory\[106\]\[6\]
+ u_cpu.rf_ram.memory\[107\]\[6\] _02005_ _01660_ _02393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_55_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10449__A1 _04562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08521_ u_cpu.rf_ram.memory\[72\]\[2\] _03647_ _03648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09303__A2 _04142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05733_ u_cpu.cpu.csr_d_sel u_cpu.cpu.decode.co_mem_word u_cpu.cpu.decode.op21 _01372_
+ _01384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_2
XFILLER_82_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06117__A2 _01724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06748__S0 _02074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08452_ _03509_ _03606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07865__A2 _03229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout39_I net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05876__A1 _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07403_ _02920_ _02921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08383_ _02845_ _03560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09067__A1 _03975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07334_ _02869_ _02870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07617__A2 _03062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07265_ _02746_ _02818_ _02821_ _00051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09004_ u_cpu.rf_ram.memory\[125\]\[4\] _03950_ _03953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06216_ u_cpu.rf_ram.memory\[132\]\[0\] u_cpu.rf_ram.memory\[133\]\[0\] u_cpu.rf_ram.memory\[134\]\[0\]
+ u_cpu.rf_ram.memory\[135\]\[0\] _01831_ _01832_ _01833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07196_ _02771_ _02772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11177__A2 _05478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06147_ u_cpu.rf_ram.memory\[92\]\[0\] u_cpu.rf_ram.memory\[93\]\[0\] u_cpu.rf_ram.memory\[94\]\[0\]
+ u_cpu.rf_ram.memory\[95\]\[0\] _01762_ _01763_ _01764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08042__A2 _03337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09790__A2 _04510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06078_ _01678_ _01695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout500 net502 net500 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_63_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout511 net515 net511 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_115_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09906_ _04611_ _04612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout522 net536 net522 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_43_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout533 net534 net533 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_104_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout544 net546 net544 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout555 net556 net555 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_86_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09837_ _04436_ _04523_ _04553_ _04554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[30\]_SI u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09768_ _04489_ _04490_ _04491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_41_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08719_ _03755_ _03766_ _03772_ _00554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09699_ _04405_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[3\] _04424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11730_ _00434_ net136 u_cpu.rf_ram.memory\[9\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_27_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07856__A2 _03215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11940__CLK net462 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11661_ _00365_ net191 u_cpu.rf_ram.memory\[19\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10612_ _05119_ _01101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07608__A2 _03049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11592_ _00296_ net245 u_cpu.rf_ram.memory\[66\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06816__B1 _02424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10543_ u_cpu.rf_ram.memory\[95\]\[4\] _05076_ _05079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08281__A2 _03495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06911__S0 _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10474_ _02787_ _05004_ _05031_ _05032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11168__A2 _05469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12213_ _00896_ net318 u_cpu.rf_ram.memory\[114\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09230__A1 _04070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12144_ _00827_ net398 u_cpu.rf_ram.memory\[115\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07792__A1 u_cpu.rf_ram.memory\[119\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_scanchain_local.scan_flop\[17\] u_arbiter.i_wb_cpu_rdt\[14\] net542 u_arbiter.i_wb_cpu_dbus_dat\[11\]
+ net11 u_arbiter.i_wb_cpu_rdt\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
X_12075_ _00758_ net318 u_cpu.rf_ram.memory\[117\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10679__A1 _05148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11026_ _05379_ _05380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_42_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11470__CLK net347 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12596__CLK net274 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06099__I _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11928_ _00624_ net333 u_cpu.rf_ram.memory\[22\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_u_scanchain_local.scan_flop\[46\]_SE net558 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05731__I u_cpu.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10851__A1 _02981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout243_I net244 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11859_ _00555_ net477 u_cpu.rf_ram.memory\[49\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout410_I net412 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08272__A2 _03488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06902__S0 _01792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07658__I _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07050_ _02647_ _02652_ _02653_ _00016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_12_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06001_ _01611_ _01617_ _01618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10084__I _04737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08024__A2 _03328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09221__A1 _04061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09772__A2 _04492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07783__A1 _03084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07952_ _03288_ _03289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__10812__I _05244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10119__B1 _04558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07393__I _02912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06903_ _01791_ _02512_ _01770_ _02513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_110_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07883_ _03179_ _03241_ _03243_ _00247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09622_ u_arbiter.i_wb_cpu_rdt\[22\] _04293_ _04359_ u_arbiter.i_wb_cpu_dbus_dat\[22\]
+ _04365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06834_ u_cpu.rf_ram.memory\[4\]\[7\] u_cpu.rf_ram.memory\[5\]\[7\] u_cpu.rf_ram.memory\[6\]\[7\]
+ u_cpu.rf_ram.memory\[7\]\[7\] _01640_ _02071_ _02444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09553_ u_arbiter.i_wb_cpu_dbus_dat\[3\] _04306_ _04311_ _04315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_110_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09288__A1 _04068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06765_ _01725_ _02375_ _02376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08504_ _03637_ _00474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05716_ _01368_ u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07838__A2 _03202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09484_ u_cpu.rf_ram.memory\[116\]\[2\] _04262_ _04263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06696_ u_cpu.rf_ram.memory\[100\]\[5\] u_cpu.rf_ram.memory\[101\]\[5\] u_cpu.rf_ram.memory\[102\]\[5\]
+ u_cpu.rf_ram.memory\[103\]\[5\] _02122_ _01895_ _02308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_58_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08435_ _03593_ _03590_ _03594_ _00448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12319__CLK net532 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06510__A2 _02123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08366_ u_cpu.rf_ram.memory\[52\]\[0\] _03550_ _03551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07317_ u_cpu.rf_ram_if.wdata0_r\[2\] u_cpu.rf_ram_if.wdata1_r\[2\] _02844_ _02857_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_123_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09460__A1 _04244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08263__A2 _03477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08297_ u_cpu.rf_ram.memory\[56\]\[6\] _03495_ _03508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06113__I2 u_cpu.rf_ram.memory\[98\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09984__S _01446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10070__A2 _04630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11343__CLK net170 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07248_ _02752_ _02806_ _02811_ _00044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08015__A2 _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07179_ _02757_ _02758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09783__I _04400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10190_ _04852_ _00946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06121__S1 _01737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11493__CLK net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout330 net332 net330 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__05816__I _01452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout341 net344 net341 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_47_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout352 net354 net352 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_28_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09515__A2 _04271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout363 net365 net363 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_82_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout374 net375 net374 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_101_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout385 net388 net385 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_87_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout396 net397 net396 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[69\]_SE net559 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09279__A1 _04056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11086__A1 _02529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11713_ _00417_ net450 u_cpu.rf_ram.memory\[53\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12693_ _01363_ net257 u_cpu.rf_ram_if.rdata0\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07679__S _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11644_ _00348_ net188 u_cpu.rf_ram.memory\[61\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09826__I0 u_arbiter.i_wb_cpu_rdt\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09987__C1 _04682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11575_ _00279_ net340 u_cpu.rf_ram.memory\[68\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06265__A1 _01691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10526_ _05053_ _05061_ _05068_ _01066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11836__CLK net487 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10457_ _05014_ _05016_ _01049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08006__A2 _03316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11010__A1 u_cpu.rf_ram.memory\[86\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09754__A2 _04477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10388_ _04972_ _04973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06407__I3 u_cpu.rf_ram.memory\[119\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06812__I0 u_cpu.rf_ram.memory\[72\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12127_ _00810_ net407 u_cpu.rf_ram.memory\[112\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10632__I _04807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12058_ _00741_ net307 u_cpu.rf_ram.memory\[35\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07517__A1 _02996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10116__A3 _04799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11009_ _05347_ _05368_ _05370_ _01247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout360_I net362 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout458_I net459 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06740__A2 _02351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11077__A1 u_cpu.rf_ram.memory\[88\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06550_ _02157_ _02159_ _02161_ _02163_ _02050_ _02164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_59_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06481_ _01638_ _02095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09690__A1 _03114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08493__A2 _03620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08220_ _03456_ _00371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11366__CLK net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08151_ u_cpu.rf_ram.memory\[61\]\[2\] _03413_ _03414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08245__A2 _03460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07388__I _02767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07102_ _02683_ _02689_ _02691_ _00022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_14_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06292__I _01652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08082_ u_cpu.rf_ram.memory\[29\]\[0\] _03370_ _03371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06351__S1 _01965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07033_ _02637_ _02631_ _02632_ _02639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_66_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11001__A1 _05363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08213__S _03451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06559__A2 _02172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08984_ u_cpu.rf_ram.memory\[126\]\[4\] _03938_ _03941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07935_ _03273_ _03278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07508__A1 _02989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09552__B _04285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07866_ _03228_ _03233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09605_ u_arbiter.i_wb_cpu_rdt\[16\] _04347_ _04344_ u_arbiter.i_wb_cpu_dbus_dat\[16\]
+ _04354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_28_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06895__C _01757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06817_ _02026_ _02418_ _02427_ _02428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_99_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07797_ _03070_ _03188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__12141__CLK net396 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09536_ _03132_ _04300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06748_ u_cpu.rf_ram.memory\[0\]\[6\] u_cpu.rf_ram.memory\[1\]\[6\] u_cpu.rf_ram.memory\[2\]\[6\]
+ u_cpu.rf_ram.memory\[3\]\[6\] _02074_ _01585_ _02359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06467__I _01596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11709__CLK net416 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09467_ _03912_ _04251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08484__A2 _03621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06679_ _02098_ _02290_ _01873_ _02291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08418_ _03583_ _00442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12291__CLK net495 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09398_ _04207_ _00799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06590__S1 _02099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11859__CLK net477 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08349_ _03491_ _03537_ _03540_ _00416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08236__A2 _03461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10043__A2 _02624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11240__A1 u_cpu.rf_ram.memory\[98\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11360_ _00064_ net68 u_cpu.rf_ram.memory\[20\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06798__A2 _02399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10311_ _04925_ _00994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_11291_ _05546_ _05547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10242_ _04880_ _00970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10173_ u_cpu.rf_ram.memory\[31\]\[4\] _04840_ _04843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout160 net164 net160 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout171 net172 net171 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_47_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout182 net183 net182 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout193 net194 net193 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_43_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08172__A1 u_cpu.rf_ram.memory\[60\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11389__CLK net182 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10806__A1 _05215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08475__A2 _03202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09688__I _01437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12676_ _01354_ net102 u_cpu.rf_ram.memory\[23\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06581__S1 _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11627_ _00331_ net177 u_cpu.rf_ram.memory\[63\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09424__A1 _04156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08227__A2 _03425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06238__A1 _01619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10034__A2 _04710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11558_ _00262_ net250 u_cpu.rf_ram.memory\[76\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07986__A1 _03268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10509_ u_cpu.rf_ram.memory\[97\]\[7\] _05040_ _05058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout206_I net207 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11489_ _00193_ net178 u_cpu.rf_ram.memory\[16\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06410__A1 _01423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06261__I1 u_cpu.rf_ram.memory\[41\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05981_ _01582_ _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12164__CLK net390 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07720_ _03119_ _03134_ _03137_ _03138_ _03139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_22_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07651_ _02723_ _03005_ _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06602_ _01862_ _02205_ _02214_ _02215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_111_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07582_ _02989_ _03036_ _03041_ _00148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_59_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10030__C _04419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09321_ u_cpu.rf_ram.memory\[120\]\[7\] _04141_ _04159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06533_ _01702_ _02147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08466__A2 _03609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09663__A1 _04249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06477__A1 _01649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout21_I net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09252_ _04072_ _04106_ _04114_ _00746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10273__A2 _04894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06464_ _01610_ _02078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06572__S1 _01585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08203_ u_cpu.rf_ram.memory\[19\]\[5\] _03443_ _03447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09183_ _03909_ _04068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09415__A1 u_cpu.rf_ram.memory\[112\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06395_ _02008_ _02009_ _02010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06229__A1 _01590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08134_ u_cpu.rf_ram.memory\[62\]\[5\] _03398_ _03402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09966__A2 _04665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06619__I3 u_cpu.rf_ram.memory\[119\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08065_ _03355_ _03360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07016_ _02605_ _02616_ _00728_ _02621_ _02622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_68_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12507__CLK net163 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08967_ _03913_ _03923_ _03930_ _00644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11289__A1 _02915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07918_ _03080_ _03266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_75_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08898_ _03881_ _03883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11531__CLK net489 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07849_ _03191_ _03216_ _03222_ _00234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06704__A2 _02315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06197__I _01813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10860_ _05269_ _05276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09519_ _03122_ _04283_ _04284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09654__A1 _04237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10791_ _05231_ _05233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11681__CLK net324 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06307__I2 u_cpu.rf_ram.memory\[86\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12530_ _01209_ net276 u_cpu.rf_ram.memory\[84\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10264__A2 _04894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09301__I _03899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_142_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12461_ _01140_ net37 u_cpu.rf_ram.memory\[104\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08209__A2 _02850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10016__A2 _04452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07957__S _03289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12037__CLK net284 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11412_ _00116_ net226 u_cpu.rf_ram.memory\[45\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12392_ _01071_ net198 u_cpu.rf_ram.memory\[95\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06315__S1 _01930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11343_ _00047_ net170 u_cpu.rf_ram.memory\[81\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11274_ _02888_ _05535_ _05537_ _01345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12187__CLK net497 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10225_ _04871_ _00962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10156_ _04830_ _04811_ _04831_ _00933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06943__A2 _02551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10087_ u_arbiter.i_wb_cpu_rdt\[17\] u_arbiter.i_wb_cpu_rdt\[1\] _01441_ _04774_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_47_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08145__A1 _03405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08448__A2 _03591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout156_I net157 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10989_ _05354_ _05349_ _05356_ _01241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_43_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06459__A1 _01958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10255__A2 _04888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12659_ _01338_ net160 u_cpu.rf_ram.memory\[100\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09948__A2 _04647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06180_ _01683_ _01797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_141_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11404__CLK net221 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09870_ _04481_ _04526_ _04585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08384__A1 _03285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11554__CLK net241 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07187__A2 _02763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09581__B1 _04331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06234__I1 u_cpu.rf_ram.memory\[21\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08821_ _03813_ _03835_ _03837_ _00591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08752_ _03745_ _03790_ _03792_ _00567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06490__S0 _01686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05964_ u_cpu.raddr\[0\] _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_61_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08136__A1 u_cpu.rf_ram.memory\[62\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout69_I net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05914__I _01451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07703_ _03122_ _03123_ _03124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_94_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08683_ _03746_ _03748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05895_ _01473_ _01522_ _01523_ u_arbiter.o_wb_cpu_adr\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08687__A2 _03748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09884__A1 _04247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06242__S0 _01640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07634_ _03075_ _03064_ _03076_ _00165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10494__A2 _05047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06793__S1 _01699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07565_ u_cpu.rf_ram.memory\[41\]\[5\] _03026_ _03030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09636__A1 u_arbiter.i_wb_cpu_dbus_dat\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08439__A2 _03590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09304_ _03902_ _04147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10246__A2 _02691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06516_ _02014_ _02129_ _02130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07496_ _02981_ _02982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09121__I _02569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09235_ _02939_ _03310_ _04104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10267__I _04893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06447_ u_cpu.rf_ram.memory\[132\]\[2\] u_cpu.rf_ram.memory\[133\]\[2\] u_cpu.rf_ram.memory\[134\]\[2\]
+ u_cpu.rf_ram.memory\[135\]\[2\] _02061_ _01832_ _02062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_10_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09166_ _03988_ _04046_ _04055_ _00718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06378_ _01702_ _01993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08117_ _03351_ _03383_ _03391_ _00333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09097_ u_cpu.rf_ram.memory\[37\]\[6\] _04007_ _04012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08611__A2 _03700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06622__A1 _01647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08048_ _03347_ _03337_ _03348_ _00307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10010_ _04500_ _04698_ _04704_ _04705_ _00913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_62_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08401__S _03561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10182__A1 _02699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09999_ u_cpu.cpu.immdec.imm30_25\[3\] _04667_ _04695_ u_cpu.cpu.immdec.imm30_25\[4\]
+ _04696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_9_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11961_ _00657_ net445 u_cpu.rf_ram.memory\[125\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10912_ _05280_ _05302_ _05309_ _01211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06689__B2 _02300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11892_ _00588_ net468 u_cpu.rf_ram.memory\[133\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06784__S1 _01576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10843_ _05211_ _05257_ _05264_ _01187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09627__A1 u_arbiter.i_wb_cpu_rdt\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10774_ u_cpu.rf_ram.memory\[105\]\[1\] _05221_ _05223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12513_ _01192_ net203 u_cpu.rf_ram.memory\[108\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11427__CLK net420 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08850__A2 _03847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07687__S _03101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12444_ _01123_ net76 u_cpu.rf_ram.memory\[102\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[47\] u_scanchain_local.module_data_in\[46\] net558 u_arbiter.o_wb_cpu_adr\[9\]
+ net26 u_scanchain_local.module_data_in\[47\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_86_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12375_ _01054_ net74 u_cpu.rf_ram.memory\[97\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08602__A2 _03698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11577__CLK net347 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06390__I _01620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11326_ _00030_ net91 u_cpu.rf_ram.memory\[82\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06323__C _01807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11257_ _05522_ _05527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07169__A2 u_cpu.rf_ram_if.wdata1_r\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10208_ _04862_ _00954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11188_ u_cpu.rf_ram.memory\[25\]\[6\] _05481_ _05486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06916__A2 _02525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10139_ u_cpu.rf_ram.memory\[32\]\[2\] _04818_ _04819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08118__A1 u_cpu.rf_ram.memory\[63\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout273_I net274 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09866__A1 _04426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08669__A2 _03734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12202__CLK net360 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout440_I net442 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout538_I net539 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07350_ _02858_ u_cpu.rf_ram.memory\[7\]\[2\] _02879_ _02882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06301_ _01761_ _01916_ _01917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07281_ _02830_ _02831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08841__A2 _03847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09020_ u_cpu.rf_ram.memory\[124\]\[2\] _03962_ _03963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06232_ _01840_ _01843_ _01845_ _01847_ _01607_ _01848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_34_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06163_ _01632_ _01780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07396__I _02777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[64\]_CLK net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06094_ _01605_ _01711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09922_ _02679_ _02703_ _01377_ _02529_ _04627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__09825__B _04542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09853_ _04470_ _04566_ _04568_ _04419_ _04569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_8_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08221__S _03450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08804_ _03824_ _03816_ _03825_ _00586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09784_ _04504_ _04505_ _04506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_74_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06996_ _02591_ _02602_ _02603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08109__A1 _03342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08735_ _03777_ _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05947_ _01406_ _01564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09857__A1 _04558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09857__B2 _04572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10467__A2 _05025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08666_ _03671_ _03734_ _03737_ _00536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05878_ u_cpu.cpu.ctrl.o_ibus_adr\[16\] _01508_ _01511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_82_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06766__S1 _02099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07617_ _03018_ _03062_ _03063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10198__S _04855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08597_ u_cpu.rf_ram.memory\[70\]\[6\] _03691_ _03696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05894__A2 _01481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07548_ _02939_ _03018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_74_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[17\]_CLK net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07096__A1 _02684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07479_ u_cpu.rf_ram.memory\[45\]\[1\] _02970_ _02972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08832__A2 _03836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09218_ u_cpu.rf_ram.memory\[92\]\[0\] _04094_ _04095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10490_ u_cpu.rf_ram.memory\[97\]\[1\] _05042_ _05045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09149_ _04044_ _04046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07399__A2 _02894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08596__A1 _03680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12160_ _00843_ net311 u_cpu.rf_ram.memory\[33\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11111_ u_cpu.cpu.decode.co_ebreak _04034_ _04031_ _02562_ _05435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_85_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09735__B _04459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12091_ _00774_ net403 u_cpu.rf_ram.memory\[118\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11042_ _05363_ _05381_ _05389_ _01261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10155__A1 u_cpu.rf_ram.memory\[32\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08899__A2 _03883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07020__A1 _02569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06454__S0 _01583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12225__CLK net359 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07571__A2 _02936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09848__A1 _04545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10458__A2 _04509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11944_ _00640_ net461 u_cpu.rf_ram.memory\[127\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06757__S1 _01625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11875_ _00571_ net519 u_cpu.rf_ram.memory\[135\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12375__CLK net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10826_ u_cpu.rf_ram.memory\[107\]\[6\] _05249_ _05254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06509__S1 _01895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07087__A1 _02673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10757_ _04823_ _05211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08823__A2 _03835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09696__I _04420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10688_ _05163_ _05168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_12_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12427_ _01106_ net364 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10635__I _05131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout119_I net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08587__A1 _03671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12358_ _01037_ net127 u_cpu.rf_ram.memory\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11309_ _02915_ _05548_ _05557_ _01360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_12289_ _00972_ net500 u_arbiter.i_wb_cpu_dbus_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout390_I net391 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09000__A2 _03950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout488_I net489 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07011__A1 _02556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07011__B2 _01411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06850_ u_cpu.rf_ram.memory\[48\]\[7\] u_cpu.rf_ram.memory\[49\]\[7\] u_cpu.rf_ram.memory\[50\]\[7\]
+ u_cpu.rf_ram.memory\[51\]\[7\] _01812_ _02092_ _02460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_99_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10697__A2 _05168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10941__I0 _04184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05801_ _01447_ _01444_ _01448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06781_ _02117_ _02391_ _02392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08520_ _03642_ _03647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10449__A2 _04700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05732_ u_cpu.cpu.decode.op21 _01381_ _01382_ _01383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__08775__I _03801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06748__S1 _01585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08451_ _03604_ _03591_ _03605_ _00453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07402_ _02721_ _02919_ _02920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_23_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08382_ _03510_ _03550_ _03559_ _00430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11742__CLK net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07078__A1 _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07333_ u_cpu.rf_ram_if.wdata0_r\[6\] u_cpu.rf_ram_if.wdata1_r\[6\] _02736_ _02869_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_17_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07264_ u_cpu.rf_ram.memory\[18\]\[1\] _02819_ _02821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07093__A4 _02682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09003_ _03907_ _03946_ _03952_ _00658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06215_ _01788_ _01832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07195_ _02734_ u_cpu.rf_ram_if.wdata0_r\[6\] _02770_ _02771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__11892__CLK net468 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06146_ _01687_ _01763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_118_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10385__A1 u_cpu.rf_ram.memory\[109\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07250__A1 _02758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06077_ u_cpu.rf_ram.memory\[44\]\[0\] u_cpu.rf_ram.memory\[45\]\[0\] u_cpu.rf_ram.memory\[46\]\[0\]
+ u_cpu.rf_ram.memory\[47\]\[0\] _01692_ _01693_ _01694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_132_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout501 net502 net501 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_82_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09378__I0 _04194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09905_ _04527_ _04489_ _04611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout512 net514 net512 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout523 net527 net523 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout534 net535 net534 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout545 net546 net545 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout556 net557 net556 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09542__A3 u_arbiter.i_wb_cpu_dbus_dat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09836_ _04552_ _04553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08886__S _03872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09767_ _04432_ _04490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06979_ u_cpu.cpu.state.o_cnt_r\[0\] _02565_ _02586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08718_ u_cpu.rf_ram.memory\[49\]\[3\] _03770_ _03772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09698_ _03114_ u_arbiter.i_wb_cpu_rdt\[5\] _04422_ _04423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07305__A2 _02724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08649_ _03673_ _03722_ _03727_ _00529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_109_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11660_ _00364_ net188 u_cpu.rf_ram.memory\[19\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10611_ u_arbiter.i_wb_cpu_rdt\[22\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[6\]
+ _05117_ _05119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_23_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11591_ _00295_ net245 u_cpu.rf_ram.memory\[66\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06816__A1 _02420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10542_ _05049_ _05072_ _05078_ _01072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06667__I1 u_cpu.rf_ram.memory\[29\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06911__S1 _01616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10473_ _02701_ _05004_ _05031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_13_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06154__B _01770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12212_ _00895_ net318 u_cpu.rf_ram.memory\[114\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07965__S _03288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10376__A1 _04817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12143_ _00826_ net396 u_cpu.rf_ram.memory\[115\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10391__S _04973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09369__I0 _04188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12074_ _00757_ net312 u_cpu.rf_ram.memory\[117\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06601__C _01733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11615__CLK net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11025_ _03061_ _05243_ _05379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10679__A2 _05152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08741__A1 _03757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07544__A2 _03011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11765__CLK net514 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11927_ _00623_ net419 u_cpu.rf_ram.memory\[22\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10300__A1 u_cpu.cpu.ctrl.o_ibus_adr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10300__B2 u_cpu.cpu.ctrl.o_ibus_adr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10851__A2 _05243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11858_ _00554_ net420 u_cpu.rf_ram.memory\[49\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10809_ _04958_ _05243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_92_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout236_I net238 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11789_ _00485_ net371 u_cpu.rf_ram.memory\[72\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06902__S1 _01793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout403_I net407 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06283__A2 _01898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07480__A1 _02897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06000_ u_cpu.rf_ram.memory\[20\]\[0\] u_cpu.rf_ram.memory\[21\]\[0\] u_cpu.rf_ram.memory\[22\]\[0\]
+ u_cpu.rf_ram.memory\[23\]\[0\] _01614_ _01616_ _01617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_115_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10367__A1 _02966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06999__B _02605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07232__A1 _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07951_ _03285_ _03287_ _03288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__10119__A1 u_cpu.cpu.immdec.imm31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06830__I1 u_cpu.rf_ram.memory\[9\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06902_ u_cpu.rf_ram.memory\[76\]\[7\] u_cpu.rf_ram.memory\[77\]\[7\] u_cpu.rf_ram.memory\[78\]\[7\]
+ u_cpu.rf_ram.memory\[79\]\[7\] _01792_ _01793_ _02512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_68_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12540__CLK net293 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07882_ u_cpu.rf_ram.memory\[74\]\[0\] _03242_ _03243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08732__A1 _03745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09621_ u_arbiter.i_wb_cpu_dbus_dat\[23\] _04352_ _04364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06833_ _01399_ _02442_ _02069_ _02443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_110_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09822__C _04532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09552_ u_arbiter.i_wb_cpu_dbus_dat\[4\] _04289_ _04285_ _04313_ _04314_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_83_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout51_I net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06764_ u_cpu.rf_ram.memory\[60\]\[6\] u_cpu.rf_ram.memory\[61\]\[6\] u_cpu.rf_ram.memory\[62\]\[6\]
+ u_cpu.rf_ram.memory\[63\]\[6\] _02095_ _01633_ _02375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_23_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09288__A2 _04129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08503_ _03568_ u_cpu.rf_ram.memory\[13\]\[3\] _03633_ _03637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12690__CLK net234 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05715_ _01367_ _01368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_37_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07299__A1 _02773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09483_ _04257_ _04262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06695_ _02004_ _02306_ _01587_ _02307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_91_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08434_ u_cpu.rf_ram.memory\[142\]\[1\] _03591_ _03594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10842__A2 _05261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08365_ _03548_ _03550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07316_ _02856_ _00067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08296_ _03506_ _03507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09460__A2 _04239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07247_ u_cpu.rf_ram.memory\[81\]\[2\] _02810_ _02811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12070__CLK net282 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07178_ _02756_ _02757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10358__A1 _02571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06129_ _01702_ _01746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07223__A1 _02746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08971__A1 _03919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07774__A2 _03172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout320 net322 net320 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_82_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout331 net332 net331 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout342 net344 net342 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout353 net354 net353 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_82_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout364 net365 net364 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_28_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11788__CLK net374 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout375 net382 net375 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__08723__A1 _03759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout386 net387 net386 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_86_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09819_ _02671_ _04396_ _04537_ _00890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout397 net399 net397 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10530__A1 _05057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05832__I _01455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09279__A2 _04129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09304__I _03902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11086__A2 _02572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11712_ _00416_ net417 u_cpu.rf_ram.memory\[53\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12692_ _01362_ net252 u_cpu.rf_ram_if.rdata1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11643_ _00347_ net189 u_cpu.rf_ram.memory\[61\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09826__I1 u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09987__C2 _04558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11574_ _00278_ net133 u_cpu.rf_ram.memory\[6\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12413__CLK net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10525_ u_cpu.rf_ram.memory\[94\]\[5\] _05064_ _05068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06265__A2 _01880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07462__A1 _02904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06896__S0 _01798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[7\]_D u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10456_ _04680_ _04500_ _05015_ _04482_ _05016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__12563__CLK net159 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11010__A2 _05369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10387_ _03870_ _03310_ _04972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__07494__I _02888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12126_ _00809_ net405 u_cpu.rf_ram.memory\[112\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06812__I1 u_cpu.rf_ram.memory\[73\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12057_ _00740_ net308 u_cpu.rf_ram.memory\[35\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[13\]_SE net544 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08714__A1 _03750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07517__A2 _02985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11008_ u_cpu.rf_ram.memory\[86\]\[0\] _05369_ _05370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10521__A1 u_cpu.rf_ram.memory\[94\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout186_I net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09214__I _02730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout353_I net354 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10824__A2 _05249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06480_ _01656_ _02093_ _01867_ _02094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09690__A2 u_arbiter.i_wb_cpu_rdt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout520_I net521 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08150_ _03406_ _03413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_u_scanchain_local.out_flop_CLKN net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09442__A2 _04230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10588__A1 _05049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07101_ _02690_ _02691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08081_ _03368_ _03370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06887__S0 _02142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07032_ _02631_ _02632_ _02637_ _02638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_127_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09817__C _04493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07205__A1 _02741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout99_I net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07756__A2 _03158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08983_ _03907_ _03934_ _03940_ _00650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09833__B _04549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07934_ _03257_ _03274_ _03277_ _00264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07508__A2 _02984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07865_ _03186_ _03229_ _03232_ _00240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09604_ u_arbiter.i_wb_cpu_dbus_dat\[17\] _04352_ _04353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08181__A2 _03431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06816_ _02420_ _02422_ _02424_ _02426_ _02050_ _02427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_56_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07796_ _03186_ _03183_ _03187_ _00216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_43_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09535_ _04285_ _04298_ _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06747_ _01958_ _02357_ _02358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06319__I0 u_cpu.rf_ram.memory\[72\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09130__A1 _04031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09466_ _04249_ _04239_ _04250_ _00824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_77_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10815__A2 _05246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06678_ u_cpu.rf_ram.memory\[56\]\[5\] u_cpu.rf_ram.memory\[57\]\[5\] u_cpu.rf_ram.memory\[58\]\[5\]
+ u_cpu.rf_ram.memory\[59\]\[5\] _01871_ _02099_ _02290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_52_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12436__CLK net160 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08417_ _03568_ u_cpu.rf_ram.memory\[15\]\[3\] _03579_ _03583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_36_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09397_ _04192_ u_cpu.rf_ram.memory\[11\]\[3\] _04203_ _04207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08348_ u_cpu.rf_ram.memory\[53\]\[1\] _03538_ _03540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09433__A2 _04227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07444__A1 _02907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11240__A2 _05515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08279_ _03493_ _03494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10310_ _01484_ _04922_ _04924_ u_cpu.cpu.ctrl.o_ibus_adr\[11\] _04925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07995__A2 _03313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06798__A3 _02408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11290_ _02789_ _02877_ _05546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08404__S _03561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09197__A1 _03111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10241_ u_arbiter.i_wb_cpu_dbus_adr\[29\] u_arbiter.i_wb_cpu_dbus_adr\[28\] _04848_
+ _04880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[36\]_SE net556 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07747__A2 _03155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10172_ _04821_ _04836_ _04842_ _00938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout150 net151 net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout161 net164 net161 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_102_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout172 net173 net172 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_130_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout183 net184 net183 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_93_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06558__I0 u_cpu.rf_ram.memory\[128\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout194 net231 net194 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_74_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08172__A2 _03428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10806__A2 _05233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12675_ _01353_ net102 u_cpu.rf_ram.memory\[23\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06393__I _01777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11626_ _00330_ net177 u_cpu.rf_ram.memory\[63\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07435__A1 _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11557_ _00261_ net249 u_cpu.rf_ram.memory\[76\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07986__A2 _03300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10508_ _04832_ _05057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_109_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11953__CLK net440 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11488_ _00192_ net105 u_cpu.rf_ram.memory\[16\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09188__A1 _04070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10439_ u_cpu.rf_ram.memory\[93\]\[6\] _04997_ _05002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout101_I net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06342__B _01588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08935__A1 _03907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07738__A2 _03146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10742__A1 _02922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12309__CLK net523 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12109_ _00792_ net128 u_cpu.rf_ram.memory\[8\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06410__A2 _02013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05980_ _01596_ _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07952__I _03288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout470_I net471 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09360__A1 _04156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07650_ _03087_ _03065_ _03088_ _00169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12459__CLK net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06601_ _02207_ _02209_ _02211_ _02213_ _01733_ _02214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__07910__A2 _03260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07581_ u_cpu.rf_ram.memory\[43\]\[2\] _03040_ _03041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05921__A1 u_cpu.cpu.ctrl.o_ibus_adr\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09320_ _03918_ _04158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09112__A1 _03980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06532_ _01766_ _02145_ _02031_ _02146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09663__A2 _04384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09251_ u_cpu.rf_ram.memory\[35\]\[6\] _04109_ _04114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11483__CLK net378 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06463_ _02067_ _02070_ _02073_ _02076_ _01607_ _02077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__06477__A2 _02090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08202_ _03417_ _03439_ _03446_ _00363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09182_ _04066_ _04058_ _04067_ _00722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout14_I net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06394_ u_cpu.rf_ram.memory\[100\]\[2\] u_cpu.rf_ram.memory\[101\]\[2\] u_cpu.rf_ram.memory\[102\]\[2\]
+ u_cpu.rf_ram.memory\[103\]\[2\] _01621_ _01895_ _02009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10039__B _04466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08133_ _03347_ _03394_ _03401_ _00339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06229__A2 _01844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[59\]_SE net562 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07977__A2 _03303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08064_ _03340_ _03356_ _03359_ _00312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10981__A1 u_cpu.rf_ram.memory\[110\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07015_ _02553_ _02620_ _02621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09179__A1 _04063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10553__I _05083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08926__A1 _03900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07729__A2 _03143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08966_ u_cpu.rf_ram.memory\[127\]\[5\] _03926_ _03930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07917_ _03264_ _03254_ _03265_ _00259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08897_ _03881_ _03882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06478__I _01659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08894__S _03871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07848_ u_cpu.rf_ram.memory\[139\]\[3\] _03220_ _03222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07779_ _03078_ _03168_ _03175_ _00211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11826__CLK net152 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09518_ _02528_ _04281_ _04282_ _04283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08693__I _03497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10790_ _05231_ _05232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09654__A2 _04384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07303__S _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07665__A1 u_cpu.rf_ram.memory\[50\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09449_ _03002_ _04224_ _04238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12460_ _01139_ net45 u_cpu.rf_ram.memory\[104\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11976__CLK net265 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11411_ _00115_ net224 u_cpu.rf_ram.memory\[45\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07417__A1 _02904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12391_ _01070_ net198 u_cpu.rf_ram.memory\[95\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09738__B _04462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11342_ _00046_ net174 u_cpu.rf_ram.memory\[81\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08090__A1 _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10972__A1 _05282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08217__I0 _02861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11273_ u_cpu.rf_ram.memory\[89\]\[0\] _05536_ _05537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10224_ u_arbiter.i_wb_cpu_dbus_adr\[21\] u_arbiter.i_wb_cpu_dbus_adr\[20\] _04867_
+ _04871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_49_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10155_ u_cpu.rf_ram.memory\[32\]\[6\] _04818_ _04831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11356__CLK net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12601__CLK net374 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10086_ _04738_ _04770_ _04771_ _04773_ _00921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_59_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09342__A1 _04158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08145__A2 _03407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10988_ u_cpu.rf_ram.memory\[110\]\[2\] _05355_ _05356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06459__A2 _02072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10638__I _04813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07656__A1 u_cpu.rf_ram.memory\[50\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06703__I0 u_cpu.rf_ram.memory\[120\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12658_ _01337_ net160 u_cpu.rf_ram.memory\[100\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11609_ _00313_ net236 u_cpu.rf_ram.memory\[64\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11204__A2 _05493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12589_ _01268_ net205 u_cpu.rf_ram.memory\[87\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10963__A1 _05273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12131__CLK net436 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06631__A2 _02239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06482__I2 u_cpu.rf_ram.memory\[62\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08908__A1 u_cpu.rf_ram.memory\[22\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08384__A2 _03020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09581__A1 u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08820_ u_cpu.rf_ram.memory\[132\]\[0\] _03836_ _03837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06234__I2 u_cpu.rf_ram.memory\[22\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06395__A1 _02008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12281__CLK net525 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05963_ _01398_ _01580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08751_ u_cpu.rf_ram.memory\[135\]\[0\] _03791_ _03792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06490__S1 _02103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11849__CLK net508 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09333__A1 u_cpu.rf_ram.memory\[118\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07702_ _02694_ _02595_ _03123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_38_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05894_ u_arbiter.i_wb_cpu_dbus_adr\[20\] _01481_ _01523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08682_ _03746_ _03747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07633_ u_cpu.rf_ram.memory\[47\]\[3\] _03072_ _03076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06242__S1 _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07564_ _02994_ _03022_ _03029_ _00142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08219__S _03451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09636__A2 _04319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11999__CLK net401 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09303_ _04145_ _04142_ _04146_ _00765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06515_ u_cpu.rf_ram.memory\[124\]\[3\] u_cpu.rf_ram.memory\[125\]\[3\] u_cpu.rf_ram.memory\[126\]\[3\]
+ u_cpu.rf_ram.memory\[127\]\[3\] _02015_ _01737_ _02129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_55_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07495_ _02829_ _02919_ _02981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_16_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06446_ _01613_ _02061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09234_ _04074_ _04094_ _04103_ _00739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09165_ u_cpu.rf_ram.memory\[91\]\[7\] _04044_ _04055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06377_ _01882_ _01991_ _01992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08116_ u_cpu.rf_ram.memory\[63\]\[6\] _03386_ _03391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08072__A1 u_cpu.rf_ram.memory\[64\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09096_ _03984_ _04004_ _04011_ _00692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08047_ u_cpu.rf_ram.memory\[65\]\[4\] _03343_ _03348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06622__A2 _02225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10706__A1 u_cpu.rf_ram.memory\[104\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09572__A1 u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08375__A2 _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09998_ _02530_ _04465_ _04665_ _04695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_77_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08949_ _03918_ _03919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_92_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11960_ _00656_ net465 u_cpu.rf_ram.memory\[125\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11131__A1 u_cpu.rf_ram.memory\[27\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10911_ u_cpu.rf_ram.memory\[84\]\[4\] _05306_ _05309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06689__A2 _02296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11891_ _00587_ net470 u_cpu.rf_ram.memory\[133\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10842_ u_cpu.rf_ram.memory\[83\]\[4\] _05261_ _05264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12004__CLK net408 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09627__A2 _04312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07638__A1 _03078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10773_ _05199_ _05220_ _05222_ _01159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12512_ _01191_ net203 u_cpu.rf_ram.memory\[108\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06310__A1 _01917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12443_ _01122_ net76 u_cpu.rf_ram.memory\[102\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11198__A1 _05449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08063__A1 u_cpu.rf_ram.memory\[64\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12374_ _01053_ net74 u_cpu.rf_ram.memory\[97\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11325_ _00029_ net101 u_cpu.rf_ram.memory\[82\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09982__I _04602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11256_ _02896_ _05523_ _05526_ _01338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09915__C _04472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08366__A2 _03550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10207_ u_arbiter.i_wb_cpu_dbus_adr\[13\] u_arbiter.i_wb_cpu_dbus_adr\[12\] _04861_
+ _04862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11187_ _05458_ _05478_ _05485_ _01310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10173__A2 _04840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10138_ _04809_ _04818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_7_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09315__A1 u_cpu.rf_ram.memory\[120\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10069_ _04490_ _04438_ _04757_ _04572_ _04758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_94_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11122__A1 _02693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09866__A2 _04561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07007__I u_cpu.cpu.decode.opcode\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout266_I net267 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05750__I _01367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05983__S0 _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09222__I _04092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout433_I net434 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06300_ u_cpu.rf_ram.memory\[92\]\[1\] u_cpu.rf_ram.memory\[93\]\[1\] u_cpu.rf_ram.memory\[94\]\[1\]
+ u_cpu.rf_ram.memory\[95\]\[1\] _01762_ _01915_ _01916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07280_ _02784_ _02829_ _02830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__06301__A1 _01761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06231_ _01597_ _01846_ _01603_ _01847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_141_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11189__A1 _05460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08054__A1 _03351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06162_ _01572_ _01779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__11521__CLK net430 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12647__CLK net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10936__A1 _05284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06514__C _01900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06065__B1 _01670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06093_ _01703_ _01708_ _01709_ _01710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_132_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10036__C _04582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09921_ _01381_ _04398_ _04626_ _00903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09554__A1 _04310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08357__A2 _03541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11671__CLK net314 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09852_ _04475_ _04567_ _04568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout81_I net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10164__A2 _04837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08803_ u_cpu.rf_ram.memory\[133\]\[3\] _03822_ _03825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09783_ _04400_ _04505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06995_ _02596_ _02601_ _02602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09841__B _04557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08734_ _03750_ _03778_ _03781_ _00560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05946_ _01563_ u_arbiter.o_wb_cpu_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12027__CLK net492 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11113__A1 _02576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09857__A2 _04559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07868__A1 _03188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05877_ u_cpu.cpu.ctrl.o_ibus_adr\[16\] _01508_ _01510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08665_ u_cpu.rf_ram.memory\[39\]\[1\] _03735_ _03737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07616_ _03061_ _03062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09609__A2 _04352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08596_ _03680_ _03688_ _03695_ _00508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06540__A1 _02150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12177__CLK net387 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07547_ _03000_ _03008_ _03017_ _00137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10475__I0 _05030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07096__A2 _02586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08293__A1 u_cpu.rf_ram.memory\[56\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07478_ _02889_ _02969_ _02971_ _00114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09217_ _04092_ _04094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06429_ _01929_ _02043_ _01932_ _02044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_108_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08045__A1 _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09148_ _04044_ _04045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10927__A1 u_cpu.rf_ram.memory\[59\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08596__A2 _03688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09079_ u_cpu.rf_ram.memory\[38\]\[7\] _03990_ _04001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11110_ u_cpu.cpu.genblk3.csr.mie_mtie _05434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_11_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12090_ _00773_ net401 u_cpu.rf_ram.memory\[118\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11041_ u_cpu.rf_ram.memory\[111\]\[6\] _05384_ _05389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08348__A2 _03538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10741__I _04807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06454__S1 _01841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09848__A2 _04563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10389__S _04973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07859__A1 _03227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11943_ _00639_ net461 u_cpu.rf_ram.memory\[127\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11874_ _00570_ net518 u_cpu.rf_ram.memory\[135\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09042__I _03902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10825_ _05213_ _05246_ _05253_ _01180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_18_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07087__A2 _02678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11544__CLK net261 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10756_ _05209_ _05201_ _05210_ _01154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07331__I0 _02867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10687_ _05135_ _05164_ _05167_ _01128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12426_ _01105_ net364 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10918__A1 _05286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12357_ _01036_ net125 u_cpu.rf_ram.memory\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11308_ u_cpu.rf_ram.memory\[23\]\[7\] _05546_ _05557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12288_ _00971_ net523 u_arbiter.i_wb_cpu_dbus_adr\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08339__A2 _03529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10651__I _04826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11239_ _05451_ _05511_ _05516_ _01331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09217__I _04092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout383_I net384 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05800_ _01446_ _01447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_95_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06780_ u_cpu.rf_ram.memory\[108\]\[6\] u_cpu.rf_ram.memory\[109\]\[6\] u_cpu.rf_ram.memory\[110\]\[6\]
+ u_cpu.rf_ram.memory\[111\]\[6\] _02001_ _01615_ _02391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_55_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09839__A2 _04551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06770__A1 _01772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05731_ u_cpu.cpu.decode.co_ebreak _01382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA_fanout550_I net551 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08450_ u_cpu.rf_ram.memory\[142\]\[6\] _03596_ _03605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07401_ _02783_ _02918_ _02919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_17_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08381_ u_cpu.rf_ram.memory\[52\]\[7\] _03548_ _03559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07332_ _02868_ _00071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07078__A2 _02660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08791__I _03815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10082__A1 _04469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07263_ _02740_ _02818_ _02820_ _00050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06676__I2 u_cpu.rf_ram.memory\[62\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06214_ _01613_ _01831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09002_ u_cpu.rf_ram.memory\[125\]\[3\] _03950_ _03952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08027__A1 _03268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07194_ _02748_ u_cpu.rf_ram_if.wdata1_r\[6\] _02770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_117_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10909__A1 u_cpu.rf_ram.memory\[84\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10047__B _04739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06145_ _01612_ _01762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06428__I2 u_cpu.rf_ram.memory\[70\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07250__A2 _02806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06076_ _01659_ _01693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09527__A1 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09904_ _04546_ _04609_ _04610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout502 net505 net502 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_28_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout513 net514 net513 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout524 net527 net524 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_82_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout535 net536 net535 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout546 net551 net546 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_8_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09835_ _04416_ _04472_ _04552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout557 net564 net557 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__07002__A2 u_cpu.cpu.ctrl.i_iscomp vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09766_ _04439_ _04489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_41_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06978_ u_cpu.cpu.alu.cmp_r _02585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_86_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08717_ _03752_ _03766_ _03771_ _00553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05929_ _01524_ _01549_ _01550_ u_arbiter.o_wb_cpu_adr\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09697_ _04405_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[5\] _04422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08648_ u_cpu.rf_ram.memory\[138\]\[2\] _03726_ _03727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11567__CLK net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06364__I1 u_cpu.rf_ram.memory\[49\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08579_ u_cpu.rf_ram.memory\[71\]\[7\] _03667_ _03685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10610_ _05118_ _01100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08266__A1 _03423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08407__S _03561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11590_ _00294_ net253 u_cpu.rf_ram.memory\[67\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10073__A1 _04652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07311__S _02852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10541_ u_cpu.rf_ram.memory\[95\]\[3\] _05076_ _05078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10472_ _04525_ _04613_ _05029_ _05030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12211_ _00894_ net353 u_cpu.cpu.decode.op22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10376__A2 _04961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10620__I0 u_arbiter.i_wb_cpu_rdt\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12142_ _00825_ net317 u_cpu.rf_ram.memory\[115\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09518__A1 _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12073_ _00756_ net310 u_cpu.rf_ram.memory\[117\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11024_ _05365_ _05369_ _05378_ _01254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06052__I0 u_cpu.rf_ram.memory\[60\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08741__A2 _03778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06752__A1 _02078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11926_ _00622_ net237 u_cpu.rf_ram.memory\[12\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[63\]_CLK net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10300__A2 _04915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09701__S _04417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11857_ _00553_ net420 u_cpu.rf_ram.memory\[49\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10808_ _05217_ _05233_ _05242_ _01174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11788_ _00484_ net374 u_cpu.rf_ram.memory\[72\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10064__A1 _04532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06807__A2 _02413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout131_I net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10739_ u_cpu.rf_ram.memory\[99\]\[7\] _05187_ _05198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08009__A1 _03270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07480__A2 _02969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12409_ _01088_ net81 u_cpu.rf_ram.memory\[28\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10611__I0 u_arbiter.i_wb_cpu_rdt\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09509__A1 _04249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07950_ _03286_ _03287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08980__A2 _03938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10119__A2 _04630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06901_ _01684_ _02510_ _02511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07881_ _03240_ _03242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_u_scanchain_local.scan_flop\[16\]_CLK net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09620_ _04363_ _00865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08732__A2 _03778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06832_ u_cpu.rf_ram.memory\[12\]\[7\] u_cpu.rf_ram.memory\[13\]\[7\] u_cpu.rf_ram.memory\[14\]\[7\]
+ u_cpu.rf_ram.memory\[15\]\[7\] _01813_ _01815_ _02442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_116_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07690__I _03111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06743__A1 _01637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09551_ _04289_ _03126_ _04313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06763_ _01569_ _02373_ _01602_ _02374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_71_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08502_ _03636_ _00473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05714_ u_cpu.rf_ram_if.rcnt\[2\] u_cpu.rf_ram_if.rcnt\[1\] _01366_ _01367_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09482_ _04242_ _04258_ _04261_ _00829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout44_I net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06694_ u_cpu.rf_ram.memory\[104\]\[5\] u_cpu.rf_ram.memory\[105\]\[5\] u_cpu.rf_ram.memory\[106\]\[5\]
+ u_cpu.rf_ram.memory\[107\]\[5\] _02005_ _01892_ _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_52_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08433_ _03490_ _03593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_75_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08364_ _03548_ _03549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06259__B1 _01870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09996__A1 _04692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07315_ _02855_ u_cpu.rf_ram.memory\[1\]\[1\] _02852_ _02856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_36_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08295_ _02771_ _03506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07246_ _02805_ _02810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09748__A1 _04404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07177_ _02735_ u_cpu.rf_ram_if.wdata0_r\[3\] _02755_ _02756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__10358__A2 _01412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10602__I0 u_arbiter.i_wb_cpu_rdt\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06128_ _01740_ _01743_ _01744_ _01745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07223__A2 _02792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12365__CLK net210 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08971__A2 _03923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06059_ _01675_ _01676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout310 net311 net310 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__11307__A1 _02912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout321 net322 net321 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout332 net335 net332 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout343 net344 net343 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_82_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout354 net355 net354 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_115_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout365 net366 net365 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout376 net381 net376 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_47_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout387 net388 net387 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
X_09818_ _04493_ _04477_ _04536_ _04395_ _04537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__08723__A2 _03767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08696__I _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout398 net399 net398 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_46_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06734__A1 _01830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09749_ _04470_ _04472_ _04473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11086__A3 _02565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11711_ _00415_ net331 u_cpu.rf_ram.memory\[53\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12691_ u_cpu.rf_ram_if.wtrig0 net342 u_cpu.rf_ram_if.genblk1.wtrig0_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06593__S0 _01686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11642_ _00346_ net189 u_cpu.rf_ram.memory\[61\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09320__I _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11573_ _00277_ net134 u_cpu.rf_ram.memory\[6\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06345__S0 _01959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10524_ _05051_ _05060_ _05067_ _01065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07462__A2 _02954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06896__S1 _01799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09739__A1 _04404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10455_ u_cpu.cpu.immdec.imm11_7\[1\] _02700_ _05004_ _05015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_13_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10386_ _04833_ _04962_ _04971_ _01023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06612__C _01900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[22\] u_arbiter.i_wb_cpu_rdt\[19\] net545 u_arbiter.i_wb_cpu_dbus_dat\[16\]
+ net13 u_arbiter.i_wb_cpu_rdt\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__08962__A2 _03926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12125_ _00808_ net406 u_cpu.rf_ram.memory\[112\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12056_ _00739_ net271 u_cpu.rf_ram.memory\[92\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11007_ _05367_ _05369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06725__A1 _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10521__A2 _05064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout179_I net183 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11909_ _00605_ net462 u_cpu.rf_ram.memory\[131\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout346_I net349 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07150__A1 _02723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06584__S0 _01863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12238__CLK net341 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10037__A1 _04729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09978__A1 _04563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout513_I net514 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07100_ _02602_ _02690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_14_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08080_ _03368_ _03369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08650__A1 u_cpu.rf_ram.memory\[138\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06887__S1 _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07031_ u_cpu.cpu.ctrl.pc_plus_offset_cy_r _02636_ _02637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__12388__CLK net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07205__A2 _02778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06264__I0 u_cpu.rf_ram.memory\[44\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08982_ u_cpu.rf_ram.memory\[126\]\[3\] _03938_ _03940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06964__A1 _02571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07933_ u_cpu.rf_ram.memory\[75\]\[1\] _03275_ _03277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07864_ u_cpu.rf_ram.memory\[77\]\[1\] _03230_ _03232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06716__A1 _02147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09603_ _04318_ _04352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06815_ _01791_ _02425_ _01770_ _02426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_83_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07795_ u_cpu.rf_ram.memory\[119\]\[1\] _03184_ _03187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06192__A2 _01785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09534_ _03125_ net36 _04286_ _04298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_3_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06746_ u_cpu.rf_ram.memory\[4\]\[6\] u_cpu.rf_ram.memory\[5\]\[6\] u_cpu.rf_ram.memory\[6\]\[6\]
+ u_cpu.rf_ram.memory\[7\]\[6\] _01959_ _02071_ _02357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_37_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06319__I1 u_cpu.rf_ram.memory\[73\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09465_ u_cpu.rf_ram.memory\[115\]\[4\] _04245_ _04250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06677_ _01725_ _02288_ _02289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06575__S0 _01849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08416_ _03582_ _00441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09396_ _04206_ _00798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10028__A1 _04487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09969__A1 _01443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11605__CLK net243 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08347_ _03485_ _03537_ _03539_ _00415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08278_ _02750_ _03493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07444__A2 _02942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07229_ u_cpu.rf_ram.memory\[21\]\[4\] _02796_ _02799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07595__I _03047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10240_ _04879_ _00969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11755__CLK net491 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10171_ u_cpu.rf_ram.memory\[31\]\[3\] _04840_ _04842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06004__I _01620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout140 net142 net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_47_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout151 net155 net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout162 net163 net162 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_102_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout173 net194 net173 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout184 net193 net184 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_74_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout195 net196 net195 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__10503__A2 _05047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06558__I1 u_cpu.rf_ram.memory\[129\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10397__S _04973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06566__S0 _01574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12674_ _00025_ net256 u_cpu.rf_ram.regzero vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11625_ _00329_ net176 u_cpu.rf_ram.memory\[63\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12530__CLK net276 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11556_ _00260_ net249 u_cpu.rf_ram.memory\[76\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07435__A2 _02942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10507_ _05055_ _05042_ _05056_ _01059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11487_ _00191_ net99 u_cpu.rf_ram.memory\[16\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09188__A2 _04059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10438_ _04827_ _04994_ _05001_ _01045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07199__A1 _02741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08935__A2 _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09934__B _04636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10369_ _04960_ _04962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06946__A1 _02553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10742__A2 _03061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12108_ _00791_ net117 u_cpu.rf_ram.memory\[8\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06410__A3 _02024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout296_I net297 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12039_ _00722_ net285 u_cpu.rf_ram.memory\[90\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09360__A2 _04174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06600_ _01993_ _02212_ _01996_ _02213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07580_ _03035_ _03040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_111_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05921__A2 _01537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10258__A1 _04888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06531_ u_cpu.rf_ram.memory\[88\]\[3\] u_cpu.rf_ram.memory\[89\]\[3\] u_cpu.rf_ram.memory\[90\]\[3\]
+ u_cpu.rf_ram.memory\[91\]\[3\] _02029_ _01768_ _02145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_94_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09250_ _04070_ _04106_ _04113_ _00745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06462_ _01597_ _02075_ _01603_ _02076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_21_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08201_ u_cpu.rf_ram.memory\[19\]\[4\] _03443_ _03446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09181_ u_cpu.rf_ram.memory\[90\]\[3\] _04064_ _04067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06393_ _01777_ _02008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08132_ u_cpu.rf_ram.memory\[62\]\[4\] _03398_ _03401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11778__CLK net152 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08505__S _03633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08063_ u_cpu.rf_ram.memory\[64\]\[1\] _03357_ _03359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07014_ _02617_ _02618_ _02620_ _00728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09179__A2 _04058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08926__A2 _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08965_ _03910_ _03922_ _03929_ _00643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07916_ u_cpu.rf_ram.memory\[76\]\[4\] _03260_ _03265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08896_ _03367_ _03287_ _03881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12403__CLK net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09351__A2 _04177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07847_ _03188_ _03216_ _03221_ _00233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08974__I _03933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07778_ u_cpu.rf_ram.memory\[40\]\[4\] _03172_ _03175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10249__A1 _02675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09517_ _01370_ _04034_ _04282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06729_ _02026_ _02331_ _02340_ _02341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_77_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06548__S0 _02047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12553__CLK net212 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06708__B _01709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09448_ _03893_ _04237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09379_ _04195_ _00792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10945__S _05326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11410_ _00114_ net224 u_cpu.rf_ram.memory\[45\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08415__S _03579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12390_ _01069_ net200 u_cpu.rf_ram.memory\[95\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07417__A2 _02925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11341_ _00045_ net174 u_cpu.rf_ram.memory\[81\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_4_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08090__A2 _03369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06720__S0 _01798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10972__A2 _05337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11272_ _05534_ _05536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_49_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10223_ _04870_ _00961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06928__A1 u_arbiter.i_wb_cpu_dbus_we vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09590__A2 _04338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10154_ _04829_ _04830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10085_ u_cpu.cpu.immdec.imm19_12_20\[5\] _04772_ _04773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12083__CLK net448 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10488__A1 _05039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07105__A1 _02693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10987_ _05348_ _05355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06703__I1 u_cpu.rf_ram.memory\[121\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10660__A1 _03286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12657_ _01336_ net80 u_cpu.rf_ram.memory\[98\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11608_ _00312_ net236 u_cpu.rf_ram.memory\[64\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12588_ _01267_ net201 u_cpu.rf_ram.memory\[87\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout211_I net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11539_ _00243_ net242 u_cpu.rf_ram.memory\[77\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10654__I _04829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout309_I net310 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06711__S0 _02142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10963__A2 _05336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06482__I3 u_cpu.rf_ram.memory\[63\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08908__A2 _03886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07967__I0 _02873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09581__A2 _04334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06395__A2 _02009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07592__A1 _03000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08750_ _03789_ _03791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05962_ _01570_ _01578_ _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09869__B1 _04581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10479__A1 _04493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07701_ _01374_ _02556_ _03122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09333__A2 _04165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08681_ _03019_ _03698_ _03746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05893_ u_cpu.cpu.ctrl.o_ibus_adr\[20\] _01519_ _01522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_93_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07344__A1 _02850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11450__CLK net334 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08392__I0 _03566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12576__CLK net168 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07632_ _03074_ _03075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_4_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07895__A2 _03245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09097__A1 u_cpu.rf_ram.memory\[37\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07563_ u_cpu.rf_ram.memory\[41\]\[4\] _03026_ _03029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xserv_1_570 io_oeb[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_94_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09302_ u_cpu.rf_ram.memory\[120\]\[1\] _04143_ _04146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06514_ _02119_ _02121_ _02124_ _02127_ _01900_ _02128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_34_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07494_ _02888_ _02980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_126_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07203__I _02777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09233_ u_cpu.rf_ram.memory\[92\]\[7\] _04092_ _04103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06445_ _01568_ _02060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09164_ _03986_ _04046_ _04054_ _00717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06376_ u_cpu.rf_ram.memory\[36\]\[2\] u_cpu.rf_ram.memory\[37\]\[2\] u_cpu.rf_ram.memory\[38\]\[2\]
+ u_cpu.rf_ram.memory\[39\]\[2\] _01698_ _01699_ _01991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_120_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08115_ _03349_ _03383_ _03390_ _00332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09095_ u_cpu.rf_ram.memory\[37\]\[5\] _04007_ _04011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08046_ _03077_ _03347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06622__A3 _02234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06473__I3 u_cpu.rf_ram.memory\[27\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09021__A1 _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10706__A2 _05177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09572__A2 _04329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09997_ _04494_ _04690_ _04693_ _04694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_27_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08948_ _02776_ _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06489__I _01687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08879_ _03871_ _03872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_3825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06769__S0 _01736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10910_ _05278_ _05302_ _05308_ _01210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11890_ _00586_ net470 u_cpu.rf_ram.memory\[133\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11943__CLK net461 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10841_ _05209_ _05257_ _05263_ _01186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06438__B _01810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10772_ u_cpu.rf_ram.memory\[105\]\[0\] _05221_ _05222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07638__A2 _03064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12511_ _01190_ net169 u_cpu.rf_ram.memory\[83\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06310__A2 _01919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12442_ _01121_ net76 u_cpu.rf_ram.memory\[102\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12373_ _01052_ net344 u_cpu.cpu.immdec.imm11_7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09260__A1 u_cpu.rf_ram.memory\[34\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11323__CLK net185 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11324_ _00028_ net174 u_cpu.rf_ram.memory\[82\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05821__A1 _01463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11255_ u_cpu.rf_ram.memory\[100\]\[1\] _05524_ _05526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09012__A1 _02981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08879__I _03871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10206_ _02690_ _04861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_45_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11186_ u_cpu.rf_ram.memory\[25\]\[5\] _05481_ _05485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06377__A2 _01991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11473__CLK net303 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10137_ _04816_ _04817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06399__I _01648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10068_ _04721_ _04751_ _04756_ _04757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_47_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[49\]_SE net558 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07877__A2 _03228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05888__A1 _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout161_I net164 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout259_I net260 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06348__B _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05983__S1 _01599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08826__A1 _03821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07629__A2 _03072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10633__A1 _02785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout426_I net429 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06152__I2 u_cpu.rf_ram.memory\[90\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06230_ u_cpu.rf_ram.memory\[0\]\[1\] u_cpu.rf_ram.memory\[1\]\[1\] u_cpu.rf_ram.memory\[2\]\[1\]
+ u_cpu.rf_ram.memory\[3\]\[1\] _01598_ _01599_ _01846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_106_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11189__A2 _05478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06161_ _01777_ _01778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08054__A2 _03338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06065__A1 _01655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06092_ _01662_ _01709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06065__B2 _01680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09920_ _04600_ _04625_ _04626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_116_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11816__CLK net477 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09003__A1 _03907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08789__I _03201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07693__I _03114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06811__B _01782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09554__A2 _04312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09851_ _04432_ _04477_ _04567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_67_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07565__A1 u_cpu.rf_ram.memory\[41\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08802_ _03497_ _03824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09782_ _04399_ _04504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06994_ _02597_ _02598_ _02600_ _02601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_fanout74_I net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08733_ u_cpu.rf_ram.memory\[136\]\[1\] _03779_ _03781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05945_ u_arbiter.i_wb_cpu_dbus_adr\[31\] _01562_ _01434_ _01563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08664_ _03666_ _03734_ _03736_ _00535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05876_ _01505_ _01506_ _01508_ _01509_ u_arbiter.o_wb_cpu_adr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__07868__A2 _03229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07615_ _02875_ _02919_ _03061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08595_ u_cpu.rf_ram.memory\[70\]\[5\] _03691_ _03695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07546_ u_cpu.rf_ram.memory\[51\]\[7\] _03006_ _03017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08817__A1 _02830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08293__A2 _03495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07477_ u_cpu.rf_ram.memory\[45\]\[0\] _02970_ _02971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09216_ _04092_ _04093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11346__CLK net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06428_ u_cpu.rf_ram.memory\[68\]\[2\] u_cpu.rf_ram.memory\[69\]\[2\] u_cpu.rf_ram.memory\[70\]\[2\]
+ u_cpu.rf_ram.memory\[71\]\[2\] _01792_ _01930_ _02043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_13_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10294__I _04906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09147_ _02731_ _03034_ _04044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08045__A2 _03337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06359_ u_cpu.rf_ram.memory\[24\]\[2\] u_cpu.rf_ram.memory\[25\]\[2\] u_cpu.rf_ram.memory\[26\]\[2\]
+ u_cpu.rf_ram.memory\[27\]\[2\] _01640_ _01642_ _01974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10927__A2 _05318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09078_ _03986_ _03992_ _04000_ _00685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11496__CLK net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05803__A1 _01432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08029_ _03270_ _03325_ _03334_ _00302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08699__I _03503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11040_ _05361_ _05381_ _05388_ _01260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07556__A1 u_cpu.rf_ram.memory\[41\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11942_ _00638_ net454 u_cpu.rf_ram.memory\[128\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07859__A2 _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05851__I _01452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11873_ _00569_ net518 u_cpu.rf_ram.memory\[135\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12121__CLK net405 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10824_ u_cpu.rf_ram.memory\[107\]\[5\] _05249_ _05253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10755_ u_cpu.rf_ram.memory\[79\]\[3\] _05207_ _05210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09481__A1 u_cpu.rf_ram.memory\[116\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12271__CLK net530 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10686_ u_cpu.rf_ram.memory\[103\]\[1\] _05165_ _05167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06685__I3 u_cpu.rf_ram.memory\[39\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12425_ _01104_ net363 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xu_scanchain_local.scan_flop\[52\] u_scanchain_local.module_data_in\[51\] net561 u_arbiter.o_wb_cpu_adr\[14\]
+ net29 u_scanchain_local.module_data_in\[52\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_103_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11839__CLK net421 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10918__A2 _05303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06047__A1 _01656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11040__A1 _05361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09784__A2 _04505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12356_ _01035_ net117 u_cpu.rf_ram.memory\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07795__A1 u_cpu.rf_ram.memory\[119\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06598__A2 _02210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11307_ _02912_ _05548_ _05556_ _01359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_141_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12287_ _00970_ net502 u_arbiter.i_wb_cpu_dbus_adr\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11989__CLK net263 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11238_ u_cpu.rf_ram.memory\[98\]\[2\] _05515_ _05516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07547__A1 _03000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11169_ _05460_ _05466_ _05474_ _01303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout376_I net381 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05730_ u_cpu.cpu.decode.op26 _01381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_76_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout543_I net546 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07400_ _02578_ _02714_ _02918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_51_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11369__CLK net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08380_ _03507_ _03550_ _03558_ _00429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12614__CLK net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07331_ _02867_ u_cpu.rf_ram.memory\[1\]\[5\] _02851_ _02868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_36_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09472__A1 _04253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10082__A2 _04760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07262_ u_cpu.rf_ram.memory\[18\]\[0\] _02819_ _02820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09001_ _03903_ _03946_ _03951_ _00657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06213_ _01568_ _01830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08027__A2 _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09224__A1 _04063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07193_ _02741_ _02768_ _02769_ _00031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06038__A1 _01649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11031__A1 _05352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09775__A2 _04493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06144_ _01648_ _01761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06428__I3 u_cpu.rf_ram.memory\[71\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06075_ _01620_ _01692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_67_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09903_ _04489_ _04432_ _04609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__09527__A2 _01450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout503 net505 net503 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout514 net515 net514 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_28_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout525 net527 net525 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout536 net537 net536 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout547 net550 net547 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09834_ _04545_ _04547_ _04550_ _04551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_63_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout558 net560 net558 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_100_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10393__I0 _04190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09765_ _04412_ _04486_ _04487_ _04488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_100_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06977_ _02559_ _02581_ _02583_ _02584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12144__CLK net398 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06761__A2 _02371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08716_ u_cpu.rf_ram.memory\[49\]\[2\] _03770_ _03771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05928_ u_arbiter.i_wb_cpu_dbus_adr\[27\] _01539_ _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09696_ _04420_ _04421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08647_ _03721_ _03726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10845__A1 _05213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05859_ _01495_ _01492_ _01496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07710__A1 _01409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06513__A2 _02126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06364__I2 u_cpu.rf_ram.memory\[50\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08578_ _03509_ _03684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_70_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07529_ _03006_ _03007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09463__A1 _04247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08266__A2 _03474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10073__A2 _04760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10540_ _05046_ _05072_ _05077_ _01071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11270__A1 _02730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10471_ _04510_ _04560_ _05028_ _04701_ _05029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08018__A2 _03328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10953__S _05325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09215__A1 _04091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12210_ _00893_ net352 u_cpu.cpu.decode.op21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__11022__A1 _05363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08423__S _03578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07777__A1 _03075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12141_ _00824_ net396 u_cpu.rf_ram.memory\[115\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12072_ _00755_ net284 u_cpu.rf_ram.memory\[34\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11023_ u_cpu.rf_ram.memory\[86\]\[7\] _05367_ _05378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06201__A1 _01400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11089__A1 _02693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11511__CLK net320 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10836__A1 _05204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11925_ _00621_ net236 u_cpu.rf_ram.memory\[12\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07701__A1 _01374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06060__S0 _01674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11856_ _00552_ net422 u_cpu.rf_ram.memory\[49\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10807_ u_cpu.rf_ram.memory\[106\]\[7\] _05231_ _05242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11787_ _00483_ net350 u_cpu.rf_ram.memory\[72\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08257__A2 _03477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11661__CLK net191 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08501__I0 _03566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11261__A1 _02903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10738_ _05146_ _05189_ _05197_ _01149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08009__A2 _03313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10669_ _05137_ _05151_ _05156_ _01121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout124_I net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09206__B2 _02589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12017__CLK net450 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12408_ _01087_ net81 u_cpu.rf_ram.memory\[28\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10611__I1 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10662__I _05150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12339_ _01019_ net165 u_cpu.rf_ram.memory\[109\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06440__A1 _01400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout493_I net494 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12167__CLK net389 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06991__A2 _01371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06900_ u_cpu.rf_ram.memory\[72\]\[7\] u_cpu.rf_ram.memory\[73\]\[7\] u_cpu.rf_ram.memory\[74\]\[7\]
+ u_cpu.rf_ram.memory\[75\]\[7\] _01762_ _01763_ _02510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_68_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07880_ _03240_ _03241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07971__I _03298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08193__A1 _03405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06831_ _01637_ _02440_ _02441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09550_ _04311_ _04312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06762_ u_cpu.rf_ram.memory\[48\]\[6\] u_cpu.rf_ram.memory\[49\]\[6\] u_cpu.rf_ram.memory\[50\]\[6\]
+ u_cpu.rf_ram.memory\[51\]\[6\] _01812_ _02092_ _02373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08501_ _03566_ u_cpu.rf_ram.memory\[13\]\[2\] _03633_ _03636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05713_ u_cpu.rf_ram_if.rcnt\[0\] _01366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10827__A1 _05215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09481_ u_cpu.rf_ram.memory\[116\]\[1\] _04259_ _04261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06693_ _02117_ _02304_ _02305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08432_ _03588_ _03590_ _03592_ _00447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout37_I net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08363_ _02831_ _03425_ _03548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09445__A1 _04156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07314_ _02854_ _02855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06259__A1 _01865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10055__A2 _04739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09996__A2 _04575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08294_ _03504_ _03488_ _03505_ _00396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10058__B _04474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06354__S1 _01968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07245_ _02746_ _02806_ _02809_ _00043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11004__A1 _05365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09748__A2 u_arbiter.i_wb_cpu_rdt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07176_ _02748_ u_cpu.rf_ram_if.wdata1_r\[3\] _02755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_30_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07759__A1 _03081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06127_ _01678_ _01744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12704__D u_cpu.cpu.o_wdata1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06058_ _01658_ _01675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout300 net304 net300 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06821__I3 u_cpu.rf_ram.memory\[143\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout311 net315 net311 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_8_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11307__A2 _05548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout322 net323 net322 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_47_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout333 net334 net333 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_115_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout344 net345 net344 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout355 net356 net355 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_43_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08184__A1 _03419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout366 net367 net366 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_82_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11534__CLK net488 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09920__A2 _04625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09817_ _04484_ _04485_ _04525_ _04535_ _04493_ _04536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
Xfanout377 net381 net377 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout388 net392 net388 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_98_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout399 net402 net399 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_28_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06734__A2 _02345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06290__S0 _01741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10118__I0 u_arbiter.i_wb_cpu_rdt\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09748_ _04404_ u_arbiter.i_wb_cpu_rdt\[1\] _04471_ _04472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_27_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09679_ _03114_ _04404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_76_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08487__A2 _03625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11684__CLK net300 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11710_ _00414_ net416 u_cpu.rf_ram.memory\[54\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12690_ u_cpu.cpu.o_wdata0 net234 u_cpu.rf_ram_if.wdata0_r\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06593__S1 _02103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11641_ _00345_ net188 u_cpu.rf_ram.memory\[61\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10747__I _04813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08239__A2 _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11243__A1 _05456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09987__A2 _04672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11572_ _00276_ net122 u_cpu.rf_ram.memory\[6\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06345__S1 _01592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10523_ u_cpu.rf_ram.memory\[94\]\[4\] _05064_ _05067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09739__A2 u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10454_ _04398_ _05011_ _05013_ _05014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_87_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10385_ u_cpu.rf_ram.memory\[109\]\[7\] _04960_ _04971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12124_ _00807_ net406 u_cpu.rf_ram.memory\[112\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06422__A1 _01778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_scanchain_local.scan_flop\[15\] u_arbiter.i_wb_cpu_rdt\[12\] net542 u_arbiter.i_wb_cpu_dbus_dat\[9\]
+ net11 u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
X_12055_ _00738_ net271 u_cpu.rf_ram.memory\[92\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08175__A1 _03410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11006_ _05367_ _05368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_81_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.input_buf_clk net1 u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08478__A2 _03622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11908_ _00604_ net461 u_cpu.rf_ram.memory\[131\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07150__A2 _02731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06584__S1 _01748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10657__I _04832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout241_I net246 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11839_ _00535_ net421 u_cpu.rf_ram.memory\[39\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout339_I net340 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11234__A1 _05444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout506_I net507 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08650__A2 _03726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07030_ u_arbiter.i_wb_cpu_ibus_adr\[0\] _02635_ _02636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06661__A1 _01786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11557__CLK net249 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06413__A1 _01761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08981_ _03903_ _03934_ _03939_ _00649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06803__I3 u_cpu.rf_ram.memory\[83\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06964__A2 u_cpu.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07932_ _03252_ _03274_ _03276_ _00263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07863_ _03179_ _03229_ _03231_ _00239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06716__A2 _02327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09602_ _04350_ _04351_ _00859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06814_ u_cpu.rf_ram.memory\[76\]\[6\] u_cpu.rf_ram.memory\[77\]\[6\] u_cpu.rf_ram.memory\[78\]\[6\]
+ u_cpu.rf_ram.memory\[79\]\[6\] _02047_ _01793_ _02425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_68_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07794_ _03067_ _03186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_84_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06192__A3 _01808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09533_ u_arbiter.i_wb_cpu_dbus_dat\[2\] _04286_ _04297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06745_ _01399_ _02355_ _02069_ _02356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_71_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08469__A2 _03613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06319__I2 u_cpu.rf_ram.memory\[74\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09464_ _03909_ _04249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10276__A2 _04898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06676_ u_cpu.rf_ram.memory\[60\]\[5\] u_cpu.rf_ram.memory\[61\]\[5\] u_cpu.rf_ram.memory\[62\]\[5\]
+ u_cpu.rf_ram.memory\[63\]\[5\] _02095_ _01633_ _02288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_52_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08415_ _03566_ u_cpu.rf_ram.memory\[15\]\[2\] _03579_ _03582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_19_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06575__S1 _01965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09395_ _04190_ u_cpu.rf_ram.memory\[11\]\[2\] _04203_ _04206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09418__A1 _04150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10028__A2 _04491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08346_ u_cpu.rf_ram.memory\[53\]\[0\] _03538_ _03539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09969__A2 u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06327__S1 _01942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12332__CLK net501 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08277_ _03491_ _03487_ _03492_ _00392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07228_ _02758_ _02792_ _02798_ _00037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07159_ _02732_ _02741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12482__CLK net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[62\]_CLK net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10170_ _04817_ _04836_ _04841_ _00937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout130 net131 net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_120_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout141 net142 net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout152 net154 net152 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__07317__S _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout163 net164 net163 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_43_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout174 net176 net174 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_43_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout185 net187 net185 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__07904__A1 _03252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout196 net202 net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_74_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06020__I _01596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07132__A2 _01414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06566__S1 _01838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12673_ _01352_ net289 u_cpu.rf_ram.memory\[89\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10019__A2 _04672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11624_ _00328_ net186 u_cpu.rf_ram.memory\[63\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[15\]_CLK net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11555_ _00259_ net242 u_cpu.rf_ram.memory\[76\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07786__I _03059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10506_ u_cpu.rf_ram.memory\[97\]\[6\] _05047_ _05056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11486_ _00190_ net376 u_cpu.raddr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10437_ u_cpu.rf_ram.memory\[93\]\[5\] _04997_ _05001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07199__A2 _02773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10368_ _04960_ _04961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06946__A2 _01391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12107_ _00790_ net118 u_cpu.rf_ram.memory\[8\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10940__I _05325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10299_ _04918_ _00989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08148__A1 _03410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08410__I _03578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12038_ _00721_ net285 u_cpu.rf_ram.memory\[90\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout191_I net192 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout289_I net290 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12205__CLK net384 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09648__A1 u_arbiter.i_wb_cpu_rdt\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout456_I net457 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09648__B2 _02547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05921__A3 _01535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06530_ _01761_ _02143_ _02144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08320__A1 _03507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06461_ u_cpu.rf_ram.memory\[0\]\[3\] u_cpu.rf_ram.memory\[1\]\[3\] u_cpu.rf_ram.memory\[2\]\[3\]
+ u_cpu.rf_ram.memory\[3\]\[3\] _02074_ _01599_ _02075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_21_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12355__CLK net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08871__A2 _03863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08200_ _03415_ _03439_ _03445_ _00362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11207__A1 _05458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09180_ _03906_ _04066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06882__A1 _01703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06392_ _02004_ _02006_ _01723_ _02007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_30_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08131_ _03345_ _03394_ _03400_ _00338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09820__A1 _04421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08062_ _03335_ _03356_ _03358_ _00311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07013_ _02618_ _02619_ _02620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10850__I _04807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08964_ u_cpu.rf_ram.memory\[127\]\[4\] _03926_ _03929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08139__A1 _03353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07915_ _03077_ _03264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08895_ _03880_ _00622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07846_ u_cpu.rf_ram.memory\[139\]\[2\] _03220_ _03221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10497__A2 _05047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07777_ _03075_ _03168_ _03174_ _00210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09516_ u_cpu.cpu.bufreg.lsb\[1\] _04034_ _04031_ _01369_ _04281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__10249__A2 _02627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06728_ _02333_ _02335_ _02337_ _02339_ _02050_ _02340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_24_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06548__S1 _01803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10297__I _04909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09447_ _04158_ _04227_ _04236_ _00819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06659_ _01958_ _02270_ _02271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08862__A2 _03860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06873__A1 _01802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09378_ _04194_ u_cpu.rf_ram.memory\[8\]\[4\] _04186_ _04195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_40_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11722__CLK net450 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08329_ _03491_ _03525_ _03528_ _00408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09811__A1 _04516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08614__A2 _03704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11340_ _00044_ net174 u_cpu.rf_ram.memory\[81\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06720__S1 _02040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11271_ _05534_ _05535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11872__CLK net511 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08378__A1 _03504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10222_ u_arbiter.i_wb_cpu_dbus_adr\[20\] u_arbiter.i_wb_cpu_dbus_adr\[19\] _04867_
+ _04870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_4_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06928__A2 _02535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10760__I _04826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10153_ _02771_ _04829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12228__CLK net360 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10084_ _04737_ _04772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09878__A1 u_cpu.rf_ram.memory\[114\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[8\] u_arbiter.i_wb_cpu_rdt\[5\] net549 u_arbiter.i_wb_cpu_dbus_dat\[2\]
+ net16 u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_43_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08550__A1 _03604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12378__CLK net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10986_ _02751_ _05354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08302__A1 _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06164__I0 u_cpu.rf_ram.memory\[84\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08853__A2 _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06864__A1 _01766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12656_ _01335_ net47 u_cpu.rf_ram.memory\[98\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11607_ _00311_ net236 u_cpu.rf_ram.memory\[64\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12587_ _01266_ net200 u_cpu.rf_ram.memory\[87\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09802__A1 _04431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08605__A2 _03701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11538_ _00242_ net234 u_cpu.rf_ram.memory\[77\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06711__S1 _01915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout204_I net208 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11469_ _00173_ net302 u_cpu.rf_ram.memory\[50\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08369__A1 _03491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09030__A2 _03957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10176__A1 _04827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09236__I _04104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07592__A2 _03037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08140__I _03059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05961_ u_cpu.rf_ram.memory\[8\]\[0\] u_cpu.rf_ram.memory\[9\]\[0\] u_cpu.rf_ram.memory\[10\]\[0\]
+ u_cpu.rf_ram.memory\[11\]\[0\] _01574_ _01577_ _01578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09869__A1 _04575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07700_ u_arbiter.i_wb_cpu_dbus_dat\[6\] _03120_ _03121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10479__A2 _04491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08680_ _03484_ _03745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_61_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05892_ _01505_ _01519_ _01520_ _01521_ u_arbiter.o_wb_cpu_adr\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_113_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08541__A1 u_cpu.rf_ram.memory\[73\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07344__A2 _02877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08392__I1 u_cpu.rf_ram.memory\[9\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07631_ _02757_ _03074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07562_ _02992_ _03022_ _03028_ _00141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_59_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09097__A2 _04007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xserv_1_571 io_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_09301_ _03899_ _04145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06513_ _01728_ _02126_ _01731_ _02127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_62_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10100__A1 _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07493_ _02916_ _02970_ _02979_ _00121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09232_ _04072_ _04094_ _04102_ _00738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06855__A1 _02098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06444_ _01947_ _02058_ _02059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_107_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09163_ u_cpu.rf_ram.memory\[91\]\[6\] _04049_ _04054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06375_ _01988_ _01989_ _01695_ _01990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_72_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08114_ u_cpu.rf_ram.memory\[63\]\[5\] _03386_ _03390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09094_ _03982_ _04003_ _04010_ _00691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08045_ _03345_ _03337_ _03346_ _00306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07280__A1 _02784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05830__A2 _01461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09021__A2 _03958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10167__A1 _04814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09996_ _04692_ _04575_ _04520_ _04693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_103_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07583__A2 _03040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08947_ _03916_ _03897_ _03917_ _00637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08878_ _03870_ _02982_ _03871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_3826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08532__A1 _03606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06769__S1 _02103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07829_ _03191_ _03204_ _03210_ _00226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06394__I0 u_cpu.rf_ram.memory\[100\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10840_ u_cpu.rf_ram.memory\[83\]\[3\] _05261_ _05263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10890__A2 _05293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12670__CLK net286 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07099__A1 _02675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10771_ _05219_ _05221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_77_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08835__A2 _03834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12510_ _01189_ net168 u_cpu.rf_ram.memory\[83\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06846__A1 _01619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12441_ _01120_ net77 u_cpu.rf_ram.memory\[102\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08599__A1 u_cpu.rf_ram.memory\[70\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12372_ _01051_ net343 u_cpu.cpu.immdec.imm11_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11323_ _00027_ net185 u_cpu.rf_ram.memory\[82\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07271__A1 u_cpu.rf_ram.memory\[18\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09399__I0 _04194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05821__A2 _01464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11254_ _02888_ _05523_ _05525_ _01337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09012__A2 _03181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10205_ _04860_ _00953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11185_ _05456_ _05477_ _05484_ _01309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10136_ _02750_ _04816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10067_ _04752_ _04726_ _04755_ _04526_ _04756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_76_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11768__CLK net481 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08523__A1 u_cpu.rf_ram.memory\[72\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05888__A2 _01516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09079__A2 _03990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10881__A2 _05290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07304__I _02845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout154_I net155 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06137__I0 u_cpu.rf_ram.memory\[116\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08826__A2 _03835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10969_ u_cpu.rf_ram.memory\[85\]\[4\] _05340_ _05343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_u_scanchain_local.scan_flop\[8\]_CLK net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06837__A1 _01786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06152__I3 u_cpu.rf_ram.memory\[91\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout321_I net322 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12639_ _01318_ net64 u_cpu.rf_ram.memory\[24\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout419_I net423 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06160_ _01397_ _01777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09251__A2 _04109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06091_ u_cpu.rf_ram.memory\[32\]\[0\] u_cpu.rf_ram.memory\[33\]\[0\] u_cpu.rf_ram.memory\[34\]\[0\]
+ u_cpu.rf_ram.memory\[35\]\[0\] _01705_ _01707_ _01708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06696__S0 _02122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05812__A2 _01453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09003__A2 _03946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12543__CLK net291 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09850_ _04565_ _04566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08801_ _03821_ _03816_ _03823_ _00585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09781_ _04502_ _04503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06993_ u_cpu.cpu.state.stage_two_req _02599_ _02600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05944_ u_cpu.cpu.ctrl.o_ibus_adr\[31\] _01561_ _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_85_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08732_ _03745_ _03778_ _03780_ _00559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_6_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout67_I net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12693__CLK net257 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08663_ u_cpu.rf_ram.memory\[39\]\[0\] _03735_ _03736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05875_ u_arbiter.i_wb_cpu_dbus_adr\[15\] _01493_ _01509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06376__I0 u_cpu.rf_ram.memory\[36\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07614_ _03059_ _03060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08594_ _03678_ _03687_ _03694_ _00507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07545_ _02998_ _03008_ _03016_ _00136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08817__A2 _03814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07476_ _02968_ _02970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09490__A2 _04262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06427_ _02039_ _02041_ _02042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09215_ _04091_ _02982_ _04092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09778__B1 _04497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09146_ _04043_ _00710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12073__CLK net310 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06358_ _01630_ _01972_ _01973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06687__S0 _01767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09077_ u_cpu.rf_ram.memory\[38\]\[6\] _03995_ _04000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06300__I0 u_cpu.rf_ram.memory\[92\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06289_ _01675_ _01905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_120_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08028_ u_cpu.rf_ram.memory\[66\]\[7\] _03323_ _03334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11910__CLK net457 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09979_ _04425_ _04566_ _04659_ _04677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_77_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10560__A1 _05046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07325__S _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11941_ _00637_ net462 u_cpu.rf_ram.memory\[128\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11872_ _00568_ net511 u_cpu.rf_ram.memory\[135\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06168__C _01784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10823_ _05211_ _05245_ _05252_ _01179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06963__I u_cpu.cpu.decode.op21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12416__CLK net357 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10754_ _04820_ _05209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_13_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10485__I _05040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10685_ _05130_ _05164_ _05166_ _01127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_12_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12424_ _01103_ net357 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[30\]_D u_arbiter.i_wb_cpu_rdt\[27\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09233__A2 _04092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06047__A2 _01661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11440__CLK net324 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[45\] u_scanchain_local.module_data_in\[44\] net559 u_arbiter.o_wb_cpu_adr\[7\]
+ net27 u_scanchain_local.module_data_in\[45\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
X_12355_ _01034_ net116 u_cpu.rf_ram.memory\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12566__CLK net162 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06678__S0 _01871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07794__I _03067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08992__A1 _02966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11306_ u_cpu.rf_ram.memory\[23\]\[6\] _05551_ _05556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12286_ _00969_ net502 u_arbiter.i_wb_cpu_dbus_adr\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06631__C _01925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11237_ _05510_ _05515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_45_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[16\]_SE net542 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11590__CLK net253 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08744__A1 u_cpu.rf_ram.memory\[136\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07547__A2 _03008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06203__I _01613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11168_ u_cpu.rf_ram.memory\[26\]\[6\] _05469_ _05474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09942__C _04520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10551__A1 _02890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10119_ u_cpu.cpu.immdec.imm31 _04630_ _04558_ _04802_ _04803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_110_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06850__S0 _01812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11099_ u_cpu.cpu.genblk3.csr.mcause3_0\[2\] _05418_ _05427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09839__A4 _04555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout271_I net275 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout369_I net372 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout536_I net537 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07330_ _02866_ _02867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12096__CLK net408 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09472__A2 _04240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07483__A1 _02900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07261_ _02817_ _02819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_73_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09000_ u_cpu.rf_ram.memory\[125\]\[2\] _03950_ _03951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06212_ _01825_ _01828_ _01829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_121_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07192_ u_cpu.rf_ram.memory\[82\]\[5\] _02753_ _02769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_u_scanchain_local.scan_flop\[21\]_D u_arbiter.i_wb_cpu_rdt\[18\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07235__A1 u_cpu.rf_ram.memory\[21\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06143_ _01565_ _01760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11031__A2 _05380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06669__S0 _01622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11220__S _05501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06822__B _01628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08983__A1 _03907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06074_ _01609_ _01691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06541__C _01925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09902_ _04402_ _04608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout504 net505 net504 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout515 net522 net515 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_98_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07538__A2 _03011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout526 net527 net526 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_101_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09833_ _04548_ _04456_ _04549_ _04550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_86_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout537 net538 net537 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout548 net549 net548 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout559 net563 net559 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10542__A1 _05049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06597__I0 u_cpu.rf_ram.memory\[36\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09764_ _04429_ _04442_ _04487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06841__S0 _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06976_ _01372_ _02581_ _02582_ _02583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05952__I _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08715_ _03765_ _03770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05927_ _01547_ _01548_ _01549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_100_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11098__A2 _01394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09695_ u_arbiter.i_wb_cpu_rdt\[6\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[6\]
+ _04417_ _04420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_26_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09160__A1 _03982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05858_ u_cpu.cpu.ctrl.o_ibus_adr\[12\] _01495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08646_ _03671_ _03722_ _03725_ _00528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12439__CLK net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07710__A2 _02559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05789_ _01436_ u_arbiter.o_wb_cpu_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08577_ _03682_ _03669_ _03683_ _00501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07528_ _03002_ _03005_ _03006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09463__A2 _04239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07474__A1 _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07459_ u_cpu.rf_ram.memory\[46\]\[2\] _02958_ _02959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11463__CLK net226 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11270__A2 _03019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10470_ _04419_ _04452_ _05025_ _04582_ _05028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA_u_scanchain_local.scan_flop\[12\]_D u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09215__A2 _02982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07226__A1 _02752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09129_ _01432_ _04032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11022__A2 _05369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[39\]_SE net552 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12140_ _00823_ net396 u_cpu.rf_ram.memory\[115\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07777__A2 _03168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05788__A1 u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12071_ _00754_ net283 u_cpu.rf_ram.memory\[34\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07119__I _02695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11022_ _05363_ _05369_ _05377_ _01253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08726__A1 u_cpu.rf_ram.memory\[49\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06023__I _01639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06201__A2 _01817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06832__S0 _01813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06052__I2 u_cpu.rf_ram.memory\[62\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11089__A2 _01393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06179__B _01795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09151__A1 _03969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11924_ _00620_ net146 u_cpu.rf_ram.memory\[12\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10836__A2 _05257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07701__A2 _02556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06060__S1 _01676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11855_ _00551_ net422 u_cpu.rf_ram.memory\[49\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11806__CLK net347 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10806_ _05215_ _05233_ _05241_ _01173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11786_ _00482_ net350 u_cpu.rf_ram.memory\[72\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06268__A2 _01883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07465__A1 u_cpu.rf_ram.memory\[46\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11261__A2 _05523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10737_ u_cpu.rf_ram.memory\[99\]\[6\] _05192_ _05197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06512__I0 u_cpu.rf_ram.memory\[96\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10668_ u_cpu.rf_ram.memory\[102\]\[2\] _05155_ _05156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12407_ _01086_ net500 u_cpu.cpu.genblk1.align.ctrl_misal vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07217__A1 _02786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11013__A2 _05372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10599_ _05112_ _01095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout117_I net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06642__B _01810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10072__I0 u_arbiter.i_wb_cpu_rdt\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08965__A1 _03910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12338_ _01018_ net167 u_cpu.rf_ram.memory\[109\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05779__A1 _01400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06361__C _01428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06440__A2 _02054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12269_ _00952_ net530 u_arbiter.i_wb_cpu_dbus_adr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08717__A1 _03752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10524__A1 _05051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06579__I0 u_cpu.rf_ram.memory\[28\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout486_I net487 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06728__B1 _02337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08193__A2 _03439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06830_ u_cpu.rf_ram.memory\[8\]\[7\] u_cpu.rf_ram.memory\[9\]\[7\] u_cpu.rf_ram.memory\[10\]\[7\]
+ u_cpu.rf_ram.memory\[11\]\[7\] _01591_ _01592_ _02440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06823__S0 _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11336__CLK net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05772__I _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07940__A2 _03278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06761_ _01697_ _02371_ _02372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09142__A1 _04032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10288__B1 _04910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08500_ _03635_ _00472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09480_ _04237_ _04258_ _04260_ _00828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06692_ u_cpu.rf_ram.memory\[108\]\[5\] u_cpu.rf_ram.memory\[109\]\[5\] u_cpu.rf_ram.memory\[110\]\[5\]
+ u_cpu.rf_ram.memory\[111\]\[5\] _02001_ _01615_ _02304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10827__A2 _05246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08431_ u_cpu.rf_ram.memory\[142\]\[0\] _03591_ _03592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11486__CLK net376 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06751__I0 u_cpu.rf_ram.memory\[20\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08362_ _03510_ _03538_ _03547_ _00422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09445__A2 _04227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07313_ u_cpu.rf_ram_if.wdata0_r\[1\] u_cpu.rf_ram_if.wdata1_r\[1\] _02844_ _02854_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06259__A2 _01868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08293_ u_cpu.rf_ram.memory\[56\]\[5\] _03495_ _03505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09996__A3 _04520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07244_ u_cpu.rf_ram.memory\[81\]\[1\] _02807_ _02809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06108__I _01665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07175_ _02733_ _02752_ _02754_ _00028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06552__B _01810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05947__I _01406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08956__A1 _03894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06126_ u_cpu.rf_ram.memory\[120\]\[0\] u_cpu.rf_ram.memory\[121\]\[0\] u_cpu.rf_ram.memory\[122\]\[0\]
+ u_cpu.rf_ram.memory\[123\]\[0\] _01741_ _01742_ _01743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07759__A2 _03155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10074__B _04553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06967__B1 _02567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06271__C _01711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06431__A2 _02045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06057_ _01673_ _01674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_47_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06282__I2 u_cpu.rf_ram.memory\[98\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout301 net303 net301 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__08708__A1 _02803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout312 net315 net312 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__06982__A3 _02546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout323 net337 net323 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_114_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout334 net335 net334 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__10515__A1 _05039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout345 net356 net345 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_113_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout356 net367 net356 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_28_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08184__A2 _03428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09816_ _04468_ _04457_ _04532_ _04534_ _04535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
Xfanout367 net394 net367 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_8_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout378 net380 net378 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__06814__S0 _02047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout389 net391 net389 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_115_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12261__CLK net491 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09154__I _04044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07931__A2 _03275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09747_ _04405_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\] _04471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_101_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10118__I1 u_arbiter.i_wb_cpu_rdt\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06959_ _02562_ _02563_ _02565_ _02566_ _02567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__06290__S1 _01905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09133__A1 _04031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08993__I _03945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10818__A2 _05249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09678_ _04399_ _04400_ _04401_ _04402_ _04403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XTAP_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07695__A1 _03115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08629_ _03715_ _00521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06727__B _01770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11640_ _00344_ net188 u_cpu.rf_ram.memory\[61\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11979__CLK net265 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09436__A2 _04230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11571_ _00275_ net114 u_cpu.rf_ram.memory\[6\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11243__A2 _05511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10451__B1 _05010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07998__A2 _03316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10522_ _05049_ _05060_ _05066_ _01064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_6_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10453_ _04560_ _05012_ _05013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10763__I _04829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06670__A2 _02281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06462__B _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08947__A1 _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10384_ _04830_ _04962_ _04970_ _01022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12123_ _00806_ net406 u_cpu.rf_ram.memory\[112\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11359__CLK net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12054_ _00737_ net270 u_cpu.rf_ram.memory\[92\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12604__CLK net378 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11005_ _05300_ _03286_ _05367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10204__S _04855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06805__S0 _01752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07922__A2 _03260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05933__A1 _01489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11907_ _00603_ net463 u_cpu.rf_ram.memory\[131\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11838_ _00534_ net478 u_cpu.rf_ram.memory\[138\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout234_I net235 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11234__A2 _05511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11769_ _00465_ net481 u_cpu.rf_ram.memory\[140\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06110__A1 _01725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12134__CLK net438 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout401_I net402 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06661__A2 _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05767__I _01417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10745__A1 u_cpu.rf_ram.memory\[79\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07610__A1 _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08980_ u_cpu.rf_ram.memory\[126\]\[2\] _03938_ _03939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12284__CLK net504 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06964__A3 _01413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07931_ u_cpu.rf_ram.memory\[75\]\[0\] _03275_ _03276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07862_ u_cpu.rf_ram.memory\[77\]\[0\] _03230_ _03231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09601_ u_arbiter.i_wb_cpu_rdt\[15\] _04347_ _04344_ u_arbiter.i_wb_cpu_dbus_dat\[15\]
+ _04351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_111_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07913__A2 _03260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06813_ _01684_ _02423_ _02424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05924__A1 _01524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07793_ _03179_ _03183_ _03185_ _00215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09115__A1 u_cpu.rf_ram.memory\[36\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09532_ _04288_ _04291_ _04296_ _00844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06744_ u_cpu.rf_ram.memory\[12\]\[6\] u_cpu.rf_ram.memory\[13\]\[6\] u_cpu.rf_ram.memory\[14\]\[6\]
+ u_cpu.rf_ram.memory\[15\]\[6\] _01813_ _01815_ _02355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_25_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09666__A2 _04388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09463_ _04247_ _04239_ _04248_ _00823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06675_ _01569_ _02286_ _01867_ _02287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06724__I0 u_cpu.rf_ram.memory\[72\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08414_ _03581_ _00440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09394_ _04205_ _00797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10069__B _04757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07429__A1 _02700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08345_ _03536_ _03538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09858__B _04573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08276_ u_cpu.rf_ram.memory\[56\]\[1\] _03488_ _03492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07227_ u_cpu.rf_ram.memory\[21\]\[3\] _02796_ _02798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06652__A2 _02264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09149__I _04044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07158_ _02739_ _02740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10736__A1 _05144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06109_ u_cpu.rf_ram.memory\[100\]\[0\] u_cpu.rf_ram.memory\[101\]\[0\] u_cpu.rf_ram.memory\[102\]\[0\]
+ u_cpu.rf_ram.memory\[103\]\[0\] _01621_ _01633_ _01726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06404__A2 _02018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07089_ _02679_ _01434_ u_arbiter.o_wb_cpu_we vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_121_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09729__I0 u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout120 net131 net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout131 net132 net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_47_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout142 net147 net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__09354__A1 _04150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout153 net154 net153 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_82_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08401__I0 _03572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout164 net173 net164 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__06168__A1 _01765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11161__A1 _05451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout175 net176 net175 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_86_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07904__A2 _03254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout186 net187 net186 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout197 net202 net197 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_101_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09106__A1 u_cpu.rf_ram.memory\[36\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07333__S _02736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07668__A1 _03084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12672_ _01351_ net288 u_cpu.rf_ram.memory\[89\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08228__I _03460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06340__A1 _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11623_ _00327_ net185 u_cpu.rf_ram.memory\[63\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06971__I _02578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08093__A1 u_cpu.rf_ram.memory\[29\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11554_ _00258_ net241 u_cpu.rf_ram.memory\[76\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06904__C _01711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10493__I _05040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10505_ _04829_ _05055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11485_ _00189_ net376 u_cpu.raddr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10436_ _04824_ _04993_ _05000_ _01044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10727__A1 _05135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08898__I _03881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10367_ _02966_ _04959_ _04960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12106_ _00789_ net125 u_cpu.rf_ram.memory\[8\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10298_ _01463_ _04915_ _04917_ u_cpu.cpu.ctrl.o_ibus_adr\[6\] _04918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08148__A2 _03407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12037_ _00720_ net284 u_cpu.rf_ram.memory\[90\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06159__A1 _01772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11152__A1 _05098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05906__A1 _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout184_I net193 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07659__A1 u_cpu.rf_ram.memory\[50\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout351_I net354 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08320__A2 _03514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06460_ _01582_ _02074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_61_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06391_ u_cpu.rf_ram.memory\[104\]\[2\] u_cpu.rf_ram.memory\[105\]\[2\] u_cpu.rf_ram.memory\[106\]\[2\]
+ u_cpu.rf_ram.memory\[107\]\[2\] _02005_ _01892_ _02006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06882__A2 _02491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08130_ u_cpu.rf_ram.memory\[62\]\[3\] _03398_ _03400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08084__A1 u_cpu.rf_ram.memory\[29\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11524__CLK net432 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10966__A1 _05275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09820__A2 _04423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08061_ u_cpu.rf_ram.memory\[64\]\[0\] _03357_ _03358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06095__B1 _01701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07831__A1 _03193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07012_ u_arbiter.i_wb_cpu_dbus_dat\[0\] u_arbiter.i_wb_cpu_dbus_dat\[8\] u_arbiter.i_wb_cpu_dbus_dat\[16\]
+ u_arbiter.i_wb_cpu_dbus_dat\[24\] u_cpu.cpu.bufreg.lsb\[0\] u_cpu.cpu.bufreg.lsb\[1\]
+ _02619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_134_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10718__A1 _05146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11674__CLK net325 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06237__I2 u_cpu.rf_ram.memory\[18\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06398__A1 _02003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout97_I net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08601__I _03201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08963_ _03907_ _03922_ _03928_ _00642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09336__A1 _04152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08139__A2 _03395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07914_ _03262_ _03254_ _03263_ _00258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08894_ _03576_ u_cpu.rf_ram.memory\[12\]\[7\] _03871_ _03880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_25_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07845_ _03215_ _03220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07898__A1 _03199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07776_ u_cpu.rf_ram.memory\[40\]\[3\] _03172_ _03174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05960__I _01576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09515_ _04255_ _04271_ _04280_ _00843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06727_ _01791_ _02338_ _01770_ _02339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10578__I _05099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08311__A2 _03517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09446_ u_cpu.rf_ram.memory\[122\]\[7\] _04225_ _04236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06322__A1 _01802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06658_ u_cpu.rf_ram.memory\[4\]\[5\] u_cpu.rf_ram.memory\[5\]\[5\] u_cpu.rf_ram.memory\[6\]\[5\]
+ u_cpu.rf_ram.memory\[7\]\[5\] _01959_ _02071_ _02270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_13_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09377_ _02863_ _04194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06873__A2 _02482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06589_ _01666_ _02201_ _02202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08075__A1 _03351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08328_ u_cpu.rf_ram.memory\[54\]\[1\] _03526_ _03528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10957__A1 _05300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07822__A1 _03179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08259_ u_cpu.rf_ram.memory\[57\]\[4\] _03477_ _03480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11270_ _02730_ _03019_ _05534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08378__A2 _03550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10221_ _04869_ _00960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10152_ _04827_ _04811_ _04828_ _00932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09327__A1 _04140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10083_ u_cpu.cpu.immdec.imm19_12_20\[6\] _04572_ _04771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06031__I _01397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08550__A2 _03656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10985_ _05352_ _05349_ _05353_ _01240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08302__A2 _03488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11547__CLK net258 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06864__A2 _02473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12655_ _01334_ net47 u_cpu.rf_ram.memory\[98\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07797__I _03070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08066__A1 u_cpu.rf_ram.memory\[64\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11606_ _00310_ net244 u_cpu.rf_ram.memory\[65\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12586_ _01265_ net205 u_cpu.rf_ram.memory\[87\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11697__CLK net452 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11537_ _00241_ net241 u_cpu.rf_ram.memory\[77\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06616__A2 _02228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06172__S0 _01787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06206__I _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11468_ _00172_ net302 u_cpu.rf_ram.memory\[50\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09945__C _04466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08369__A2 _03549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10419_ _04198_ u_cpu.rf_ram.memory\[2\]\[6\] _04982_ _04990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10176__A2 _04837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11399_ _00103_ net293 u_cpu.rf_ram.memory\[42\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06650__B _01644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout399_I net402 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09961__B _04615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05960_ _01576_ _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11125__A1 _05098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09869__A2 _04580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05891_ u_arbiter.i_wb_cpu_dbus_adr\[19\] _01512_ _01521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12322__CLK net532 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08541__A2 _03659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07630_ _03071_ _03064_ _03073_ _00164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05780__I _01401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06552__A1 _02141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07561_ u_cpu.rf_ram.memory\[41\]\[3\] _03026_ _03028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06097__B _01713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xserv_1_572 io_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_09300_ _04140_ _04142_ _04144_ _00764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06512_ u_cpu.rf_ram.memory\[96\]\[3\] u_cpu.rf_ram.memory\[97\]\[3\] u_cpu.rf_ram.memory\[98\]\[3\]
+ u_cpu.rf_ram.memory\[99\]\[3\] _02125_ _01641_ _02126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_62_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07492_ u_cpu.rf_ram.memory\[45\]\[7\] _02968_ _02979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_u_scanchain_local.scan_flop\[61\]_CLK net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10100__A2 _04700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07352__I0 _02861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12472__CLK net241 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09231_ u_cpu.rf_ram.memory\[92\]\[6\] _04097_ _04102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06443_ u_cpu.rf_ram.memory\[128\]\[2\] u_cpu.rf_ram.memory\[129\]\[2\] u_cpu.rf_ram.memory\[130\]\[2\]
+ u_cpu.rf_ram.memory\[131\]\[2\] _01826_ _01827_ _02058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_72_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout12_I net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08057__A1 _03353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09162_ _03984_ _04046_ _04053_ _00716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06374_ u_cpu.rf_ram.memory\[44\]\[2\] u_cpu.rf_ram.memory\[45\]\[2\] u_cpu.rf_ram.memory\[46\]\[2\]
+ u_cpu.rf_ram.memory\[47\]\[2\] _01692_ _01879_ _01989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_21_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08113_ _03347_ _03382_ _03389_ _00331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06607__A2 _02219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09093_ u_cpu.rf_ram.memory\[37\]\[4\] _04007_ _04010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10066__C _04474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08044_ u_cpu.rf_ram.memory\[65\]\[3\] _03343_ _03346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06116__I _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09557__A1 _03132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05955__I _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10167__A2 _04836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10411__I0 _04190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09427__I _03180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09995_ _03115_ u_arbiter.i_wb_cpu_rdt\[9\] _04691_ _04692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06091__I0 u_cpu.rf_ram.memory\[32\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08780__A2 _03806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08946_ u_cpu.rf_ram.memory\[128\]\[6\] _03904_ _03917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[14\]_CLK net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08877_ _02849_ _03870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_84_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08532__A2 _03644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07828_ u_cpu.rf_ram.memory\[129\]\[3\] _03208_ _03210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06719__C _01925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07759_ _03081_ _03155_ _03162_ _00204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07099__A2 _02627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[29\]_CLK net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10770_ _05219_ _05220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_73_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09429_ _04225_ _04226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06846__A2 _02455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08048__A1 _03347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12440_ _01119_ net77 u_cpu.rf_ram.memory\[102\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12371_ _01050_ net343 u_cpu.cpu.immdec.imm11_7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11322_ _00026_ net185 u_cpu.rf_ram.memory\[82\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07271__A2 _02822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10771__I _05219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11253_ u_cpu.rf_ram.memory\[100\]\[0\] _05524_ _05525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10204_ u_arbiter.i_wb_cpu_dbus_adr\[12\] u_arbiter.i_wb_cpu_dbus_adr\[11\] _04855_
+ _04860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07023__A2 _02624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11184_ u_cpu.rf_ram.memory\[25\]\[4\] _05481_ _05484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12345__CLK net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10135_ _04814_ _04810_ _04815_ _00928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08771__A2 _03803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10066_ _04721_ _04710_ _04753_ _04754_ _04474_ _04755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_85_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09720__A1 _04443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08523__A2 _03647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10968_ _05278_ _05336_ _05342_ _01234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06137__I1 u_cpu.rf_ram.memory\[117\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06837__A2 _02446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout147_I net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10899_ _05300_ _02831_ _05301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12638_ _01317_ net63 u_cpu.rf_ram.memory\[24\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout314_I net315 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12569_ _01248_ net204 u_cpu.rf_ram.memory\[86\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06090_ _01706_ _01707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07262__A2 _02819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06696__S1 _01895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09539__A1 u_arbiter.i_wb_cpu_rdt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08800_ u_cpu.rf_ram.memory\[133\]\[2\] _03822_ _03823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08762__A2 _03794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09780_ _04433_ _04476_ _04502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06992_ u_arbiter.i_wb_cpu_dbus_dat\[5\] _01408_ _02599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11712__CLK net417 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08731_ u_cpu.rf_ram.memory\[136\]\[0\] _03779_ _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05943_ _01560_ _01557_ _01561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11218__S _05501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08662_ _03733_ _03735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05874_ u_cpu.cpu.ctrl.o_ibus_adr\[13\] u_cpu.cpu.ctrl.o_ibus_adr\[12\] _01492_ _01507_
+ _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_82_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06376__I1 u_cpu.rf_ram.memory\[37\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07613_ _02739_ _03059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08593_ u_cpu.rf_ram.memory\[70\]\[4\] _03691_ _03694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11862__CLK net420 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07544_ u_cpu.rf_ram.memory\[51\]\[6\] _03011_ _03016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07325__I0 u_cpu.rf_ram_if.wdata0_r\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10856__I _04813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06828__A2 _02438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07475_ _02968_ _02969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09214_ _02730_ _04091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06426_ u_cpu.rf_ram.memory\[64\]\[2\] u_cpu.rf_ram.memory\[65\]\[2\] u_cpu.rf_ram.memory\[66\]\[2\]
+ u_cpu.rf_ram.memory\[67\]\[2\] _01787_ _02040_ _02041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_33_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10077__B _04602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09778__A1 _02675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09145_ _01432_ u_cpu.cpu.state.o_cnt_r\[2\] _04043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_124_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09778__B2 _04500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06357_ u_cpu.rf_ram.memory\[28\]\[2\] u_cpu.rf_ram.memory\[29\]\[2\] u_cpu.rf_ram.memory\[30\]\[2\]
+ u_cpu.rf_ram.memory\[31\]\[2\] _01631_ _01634_ _01972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_108_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06288_ _01671_ _01904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07253__A2 _02810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09076_ _03984_ _03992_ _03999_ _00684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12368__CLK net210 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08027_ _03268_ _03325_ _03333_ _00301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06439__S1 _01942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08202__A1 _03417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09950__A1 _04650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08753__A2 _03791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09950__B2 _04420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09978_ _04563_ _04661_ _04676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11392__CLK net221 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08929_ _03895_ _03904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_58_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11940_ _00636_ net462 u_cpu.rf_ram.memory\[128\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07405__I _02922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11871_ _00567_ net511 u_cpu.rf_ram.memory\[135\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10822_ u_cpu.rf_ram.memory\[107\]\[4\] _05249_ _05252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08269__A1 _03380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10076__A1 _04420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10766__I _04832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10753_ _05206_ _05201_ _05208_ _01153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10684_ u_cpu.rf_ram.memory\[103\]\[0\] _05165_ _05166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12423_ _01102_ net357 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10379__A2 _04965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12354_ _01033_ net117 u_cpu.rf_ram.memory\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07244__A2 _02807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06678__S1 _02099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11305_ _02909_ _05548_ _05555_ _01358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08992__A2 _03181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12285_ _00968_ net505 u_arbiter.i_wb_cpu_dbus_adr\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10207__S _04861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[38\] u_scanchain_local.module_data_in\[37\] net552 u_arbiter.o_wb_cpu_adr\[0\]
+ net20 u_scanchain_local.module_data_in\[38\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_5_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11236_ _05449_ _05511_ _05514_ _01330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10000__A1 _04500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09941__A1 _04505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08744__A2 _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11167_ _05458_ _05466_ _05473_ _01302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10118_ u_arbiter.i_wb_cpu_rdt\[31\] u_arbiter.i_wb_cpu_rdt\[15\] _01447_ _04802_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_23_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10450__B _04560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11098_ u_cpu.cpu.genblk3.csr.mcause3_0\[3\] _01394_ _02693_ _02684_ _05426_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_83_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06850__S1 _02092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11885__CLK net468 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10049_ u_cpu.cpu.immdec.imm19_12_20\[1\] _04741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_36_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout264_I net265 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09530__I _04294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout431_I net433 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout529_I net530 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06375__B _01695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06366__S0 _01639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08146__I _03067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07260_ _02817_ _02818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07483__A2 _02969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06211_ u_cpu.rf_ram.memory\[128\]\[0\] u_cpu.rf_ram.memory\[129\]\[0\] u_cpu.rf_ram.memory\[130\]\[0\]
+ u_cpu.rf_ram.memory\[131\]\[0\] _01826_ _01827_ _01828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07191_ _02767_ _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12510__CLK net168 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06142_ _01423_ _01734_ _01758_ _01759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__08432__A1 _03588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07235__A2 _02791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06669__S1 _01625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08983__A2 _03934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06073_ _01684_ _01689_ _01690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09901_ _04601_ _04603_ _04606_ _04607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12660__CLK net159 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout505 net506 net505 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_82_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout516 net520 net516 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_09832_ _04527_ _04549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout527 net535 net527 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout538 net539 net538 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_140_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout549 net550 net549 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10542__A2 _05072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09763_ _04472_ _04486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06975_ u_cpu.cpu.alu.i_rs1 _02547_ _01408_ _02582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_6_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06841__S1 _01599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08714_ _03750_ _03766_ _03769_ _00552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05926_ u_cpu.cpu.ctrl.o_ibus_adr\[26\] u_cpu.cpu.ctrl.o_ibus_adr\[25\] u_cpu.cpu.ctrl.o_ibus_adr\[24\]
+ _01535_ _01548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_09694_ _04418_ _04419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08645_ u_cpu.rf_ram.memory\[138\]\[1\] _03723_ _03725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05857_ _01489_ _01490_ _01492_ _01494_ u_arbiter.o_wb_cpu_adr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_26_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08576_ u_cpu.rf_ram.memory\[71\]\[6\] _03674_ _03683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12040__CLK net285 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05788_ u_arbiter.i_wb_cpu_ibus_adr\[1\] _01433_ _01436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10058__A1 _04692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07527_ _03004_ _03005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11608__CLK net236 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06357__S0 _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07474__A2 _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07458_ _02953_ _02958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08671__A1 _03676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12190__CLK net498 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06409_ _02017_ _02019_ _02021_ _02023_ _01757_ _02024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_41_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06109__S0 _01621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07389_ _02909_ _02910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09128_ u_cpu.cpu.mem_bytecnt\[0\] _04031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11758__CLK net512 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07226__A2 _02792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09059_ u_cpu.rf_ram.memory\[123\]\[7\] _03971_ _03989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05788__A2 _01433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06985__A1 _01385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10781__A2 _05224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12070_ _00753_ net282 u_cpu.rf_ram.memory\[34\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11021_ u_cpu.rf_ram.memory\[86\]\[6\] _05372_ _05377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_u_scanchain_local.scan_flop\[7\]_CLK net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06832__S1 _01815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11923_ _00619_ net153 u_cpu.rf_ram.memory\[12\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07162__A1 _02736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11854_ _00550_ net510 u_cpu.rf_ram.memory\[137\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10805_ u_cpu.rf_ram.memory\[106\]\[6\] _05236_ _05241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11785_ _00481_ net350 u_cpu.rf_ram.memory\[72\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12533__CLK net276 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10736_ _05144_ _05189_ _05196_ _01148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10667_ _05150_ _05155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12406_ _01085_ net383 u_cpu.cpu.bufreg.i_sh_signed vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10598_ u_arbiter.i_wb_cpu_rdt\[16\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[0\]
+ _05111_ _05112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_126_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10072__I1 u_arbiter.i_wb_cpu_rdt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08965__A2 _03922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12337_ _01017_ net167 u_cpu.rf_ram.memory\[109\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06976__A1 _01372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06520__S0 _02133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10772__A2 _05221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06214__I _01613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08630__S _03712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12268_ _00951_ net521 u_arbiter.i_wb_cpu_dbus_adr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11219_ _05504_ _01323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12199_ _00882_ net398 u_cpu.rf_ram.memory\[113\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10524__A2 _05060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06579__I1 u_cpu.rf_ram.memory\[29\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09525__I _03132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout381_I net382 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06823__S1 _01616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout479_I net483 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06760_ u_cpu.rf_ram.memory\[52\]\[6\] u_cpu.rf_ram.memory\[53\]\[6\] u_cpu.rf_ram.memory\[54\]\[6\]
+ u_cpu.rf_ram.memory\[55\]\[6\] _01747_ _01748_ _02371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_110_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10288__A1 u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06691_ _01760_ _02274_ _02283_ _02302_ _02303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_110_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06200__I0 u_cpu.rf_ram.memory\[136\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08430_ _03589_ _03591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_63_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08361_ u_cpu.rf_ram.memory\[53\]\[7\] _03536_ _03547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06339__S0 _01574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07312_ _02853_ _00066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08653__A1 _03678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08292_ _03503_ _03504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11900__CLK net468 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10460__A1 _04401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07243_ _02740_ _02806_ _02808_ _00042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07174_ u_cpu.rf_ram.memory\[82\]\[2\] _02753_ _02754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06267__I0 u_cpu.rf_ram.memory\[36\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08956__A2 _03922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06125_ _01675_ _01742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06967__A1 _02561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10074__C _04609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06967__B2 u_cpu.cpu.genblk3.csr.mstatus_mie vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06124__I _01673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06056_ _01571_ _01673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_47_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout302 net303 net302 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__09905__A1 _04527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08708__A2 _03380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout313 net314 net313 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout324 net325 net324 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_141_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10515__A2 _05060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout335 net336 net335 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout346 net349 net346 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__09435__I _04225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout357 net366 net357 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_09815_ _04505_ _04514_ _04533_ _04534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__12406__CLK net383 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout368 net372 net368 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__06814__S1 _01793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout379 net380 net379 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_41_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09746_ _04437_ _04470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06958_ u_cpu.cpu.decode.op26 _01413_ _02566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10279__A1 _04833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05909_ _01529_ _01534_ _01535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09677_ u_arbiter.i_wb_cpu_rdt\[7\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[7\]
+ _01438_ _04402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11430__CLK net370 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06889_ u_cpu.rf_ram.memory\[88\]\[7\] u_cpu.rf_ram.memory\[89\]\[7\] u_cpu.rf_ram.memory\[90\]\[7\]
+ u_cpu.rf_ram.memory\[91\]\[7\] _01741_ _01742_ _02499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12556__CLK net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08628_ _03566_ u_cpu.rf_ram.memory\[14\]\[2\] _03712_ _03715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07695__A2 u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09170__I _04057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[0\]_SE net552 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08559_ _03490_ _03671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11580__CLK net340 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08644__A1 _03666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07447__A2 _02946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11570_ _00274_ net60 u_cpu.rf_ram.memory\[6\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10451__A1 _04407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10521_ u_cpu.rf_ram.memory\[94\]\[3\] _05064_ _05066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10451__B2 _04469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10452_ _04468_ _04510_ _04652_ _04680_ _05012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_100_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08947__A2 _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10383_ u_cpu.rf_ram.memory\[109\]\[6\] _04965_ _04970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12122_ _00805_ net406 u_cpu.rf_ram.memory\[112\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06034__I _01650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09773__C _04495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12053_ _00736_ net270 u_cpu.rf_ram.memory\[92\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10506__A2 _05047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11004_ _05365_ _05350_ _05366_ _01246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_46_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06805__S1 _02151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07383__A1 _02904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06430__I0 u_cpu.rf_ram.memory\[72\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11906_ _00602_ net471 u_cpu.rf_ram.memory\[131\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10220__S _04867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11837_ _00533_ net487 u_cpu.rf_ram.memory\[138\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10690__A1 _05137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06209__I _01613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11768_ _00464_ net481 u_cpu.rf_ram.memory\[140\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10442__A1 _04833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10719_ u_cpu.rf_ram.memory\[104\]\[7\] _05175_ _05186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_fanout227_I net228 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11699_ _00403_ net427 u_cpu.rf_ram.memory\[55\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06653__B _02265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08938__A2 _03904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09060__A1 _03988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12429__CLK net363 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07610__A2 _03049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06264__I3 u_cpu.rf_ram.memory\[47\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07930_ _03273_ _03275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05783__I net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07861_ _03228_ _03230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_60_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07374__A1 _02897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11453__CLK net334 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09600_ u_arbiter.i_wb_cpu_dbus_dat\[16\] _04338_ _04350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11170__A2 _05464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06812_ u_cpu.rf_ram.memory\[72\]\[6\] u_cpu.rf_ram.memory\[73\]\[6\] u_cpu.rf_ram.memory\[74\]\[6\]
+ u_cpu.rf_ram.memory\[75\]\[6\] _01762_ _01763_ _02423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06421__I0 u_cpu.rf_ram.memory\[84\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07792_ u_cpu.rf_ram.memory\[119\]\[0\] _03184_ _03185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09531_ u_arbiter.i_wb_cpu_rdt\[0\] _04293_ _04295_ _03125_ _04296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09115__A2 _04019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06743_ _01637_ _02353_ _02354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07126__A1 _01387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11226__S _05500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05732__B _01382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09462_ u_cpu.rf_ram.memory\[115\]\[3\] _04245_ _04248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06674_ u_cpu.rf_ram.memory\[48\]\[5\] u_cpu.rf_ram.memory\[49\]\[5\] u_cpu.rf_ram.memory\[50\]\[5\]
+ u_cpu.rf_ram.memory\[51\]\[5\] _01812_ _02092_ _02286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_25_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout42_I net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08874__A1 _03830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06724__I1 u_cpu.rf_ram.memory\[73\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08413_ _03564_ u_cpu.rf_ram.memory\[15\]\[1\] _03579_ _03581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_91_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10681__A1 _02876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09393_ _04188_ u_cpu.rf_ram.memory\[11\]\[1\] _04203_ _04205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_36_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10069__C _04572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08344_ _03536_ _03537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06119__I _01685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09674__I0 u_arbiter.i_wb_cpu_rdt\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09823__B1 _04525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08275_ _03490_ _03491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05958__I u_cpu.raddr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07226_ _02752_ _02792_ _02797_ _00036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09051__A1 _03982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07157_ _02738_ _02739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09366__S _04186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06108_ _01665_ _01725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_65_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07088_ _02633_ _02679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_79_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07601__A2 _03052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06039_ _01595_ _01656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout110 net113 net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout121 net124 net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout132 net157 net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout143 net145 net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_82_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09354__A2 _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout154 net155 net154 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_75_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout165 net167 net165 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__06168__A2 _01771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06799__S0 _02142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout176 net184 net176 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_47_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06412__I0 u_cpu.rf_ram.memory\[92\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout187 net192 net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout198 net199 net198 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__05915__A2 _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11946__CLK net444 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09729_ u_arbiter.i_wb_cpu_rdt\[8\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[8\]
+ _01439_ _04454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06738__B _01644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10672__A1 u_cpu.rf_ram.memory\[102\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12671_ _01350_ net288 u_cpu.rf_ram.memory\[89\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06340__A2 _01954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11622_ _00326_ net174 u_cpu.rf_ram.memory\[29\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08617__A1 _03680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11553_ _00257_ net241 u_cpu.rf_ram.memory\[76\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09290__A1 _04070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10504_ _05053_ _05042_ _05054_ _01058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11326__CLK net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11484_ _00188_ net378 u_cpu.rf_ram_if.rcnt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11224__I0 _02866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10435_ u_cpu.rf_ram.memory\[93\]\[4\] _04997_ _05000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10366_ _04958_ _04959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_48_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[20\] u_arbiter.i_wb_cpu_rdt\[17\] net541 u_arbiter.i_wb_cpu_dbus_dat\[14\]
+ net9 u_arbiter.i_wb_cpu_rdt\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
X_12105_ _00788_ net125 u_cpu.rf_ram.memory\[8\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10215__S _04861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10297_ _04909_ _04917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12036_ _00719_ net284 u_cpu.rf_ram.memory\[90\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06159__A2 _01775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11152__A2 _02938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout177_I net184 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08856__A1 _03832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10663__A1 u_cpu.rf_ram.memory\[102\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout344_I net345 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08608__A1 _03671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06390_ _01620_ _02005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_33_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout511_I net515 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09281__A1 _04061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08084__A2 _03370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10966__A2 _05336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06095__A1 _01690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08060_ _03355_ _03357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06095__B2 _01710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12251__CLK net274 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09569__C1 _04327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07011_ _02556_ u_cpu.cpu.mem_bytecnt\[1\] u_cpu.cpu.mem_bytecnt\[0\] _01411_ _02618_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_66_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10718__A2 _05177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09584__A2 _04338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06237__I3 u_cpu.rf_ram.memory\[19\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08962_ u_cpu.rf_ram.memory\[127\]\[3\] _03926_ _03928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07913_ u_cpu.rf_ram.memory\[76\]\[3\] _03260_ _03263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11969__CLK net446 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09336__A2 _04161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08893_ _03879_ _00621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08395__I0 _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07844_ _03186_ _03216_ _03219_ _00232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07898__A2 _03242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10859__I _04816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07775_ _03071_ _03168_ _03173_ _00209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_77_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09514_ u_cpu.rf_ram.memory\[33\]\[7\] _04269_ _04280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06726_ u_cpu.rf_ram.memory\[76\]\[5\] u_cpu.rf_ram.memory\[77\]\[5\] u_cpu.rf_ram.memory\[78\]\[5\]
+ u_cpu.rf_ram.memory\[79\]\[5\] _02047_ _01793_ _02338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_37_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09895__I0 u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09445_ _04156_ _04227_ _04235_ _00818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06657_ _01399_ _02268_ _02069_ _02269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11349__CLK net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09376_ _04193_ _00791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06588_ u_cpu.rf_ram.memory\[60\]\[4\] u_cpu.rf_ram.memory\[61\]\[4\] u_cpu.rf_ram.memory\[62\]\[4\]
+ u_cpu.rf_ram.memory\[63\]\[4\] _02095_ _01668_ _02201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_90_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08327_ _03485_ _03525_ _03527_ _00407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09272__A1 _04072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06705__S0 _02133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10957__A2 _02786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08258_ _03415_ _03473_ _03479_ _00386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07209_ _02708_ _02710_ _02783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_10_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09024__A1 u_cpu.rf_ram.memory\[124\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06881__I0 u_cpu.rf_ram.memory\[112\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08999__I _03945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08189_ _03367_ _03310_ _03438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10220_ u_arbiter.i_wb_cpu_dbus_adr\[19\] u_arbiter.i_wb_cpu_dbus_adr\[18\] _04867_
+ _04869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07586__A1 _02994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10151_ u_cpu.rf_ram.memory\[32\]\[5\] _04818_ _04828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09327__A2 _04161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10082_ _04469_ _04760_ _04769_ _04466_ _04770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_94_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08386__I0 _03560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07889__A2 _03245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10893__A1 _05282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12124__CLK net406 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10984_ u_cpu.rf_ram.memory\[110\]\[1\] _05350_ _05353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06164__I2 u_cpu.rf_ram.memory\[86\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12654_ _01333_ net93 u_cpu.rf_ram.memory\[98\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12274__CLK net533 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11605_ _00309_ net243 u_cpu.rf_ram.memory\[65\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06915__C _01405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[68\] u_scanchain_local.module_data_in\[67\] net559 u_arbiter.o_wb_cpu_adr\[30\]
+ net27 u_scanchain_local.module_data_in\[68\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
X_12585_ _01264_ net207 u_cpu.rf_ram.memory\[87\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11536_ _00240_ net250 u_cpu.rf_ram.memory\[77\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05824__A1 _01463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06172__S1 _01788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11467_ _00171_ net301 u_cpu.rf_ram.memory\[50\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10418_ _04989_ _01037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08702__I _03506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11398_ _00102_ net301 u_cpu.rf_ram.memory\[42\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07577__A1 _02980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12371__D _01050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10349_ _04947_ _01010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07318__I _02857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06222__I _01576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout294_I net298 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11125__A2 _03033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12019_ _00702_ net428 u_cpu.rf_ram.memory\[36\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05890_ u_cpu.cpu.ctrl.o_ibus_adr\[19\] _01516_ _01520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_78_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06001__A1 _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout461_I net467 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10884__A1 _05273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout559_I net563 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07560_ _02989_ _03022_ _03027_ _00140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_59_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08149__I _03070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12617__CLK net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06511_ _01673_ _02125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_62_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xserv_1_573 io_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_22_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07491_ _02913_ _02970_ _02978_ _00120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07501__A1 _02980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09230_ _04070_ _04094_ _04101_ _00737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06442_ _01819_ _02056_ _01823_ _02057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10239__I1 u_arbiter.i_wb_cpu_dbus_adr\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09161_ u_cpu.rf_ram.memory\[91\]\[5\] _04049_ _04053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08057__A2 _03338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09254__A1 _04074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06373_ _01609_ _01988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11641__CLK net188 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10939__A2 _02938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08112_ u_cpu.rf_ram.memory\[63\]\[4\] _03386_ _03389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11061__A1 u_cpu.rf_ram.memory\[87\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09092_ _03980_ _04003_ _04009_ _00690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08043_ _03074_ _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06863__I0 u_cpu.rf_ram.memory\[32\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09557__A2 _04284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11791__CLK net373 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07568__A1 _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09994_ _01440_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[9\] _04691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_66_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10082__C _04466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06240__A1 _01630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08945_ _03915_ _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11116__A2 _01378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08876_ _03832_ _03860_ _03869_ _00614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10324__B1 _04931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05971__I _01587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07827_ _03188_ _03204_ _03209_ _00225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06543__A2 _02156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06394__I2 u_cpu.rf_ram.memory\[102\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07758_ u_cpu.rf_ram.memory\[17\]\[5\] _03158_ _03162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06709_ _02314_ _02316_ _02318_ _02320_ _02139_ _02321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_44_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07689_ net2 _03111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09493__A1 _04253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09428_ _02937_ _04224_ _04225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09359_ u_cpu.rf_ram.memory\[121\]\[6\] _04177_ _04182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08048__A2 _03337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11213__I _05500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12370_ _01049_ net359 u_cpu.cpu.immdec.imm11_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11321_ _03134_ _05564_ _01365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06854__I0 u_cpu.rf_ram.memory\[56\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07339__S _02851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11252_ _05522_ _05524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07559__A1 u_cpu.rf_ram.memory\[41\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10203_ _04859_ _00952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11183_ _05454_ _05477_ _05483_ _01308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07138__I _02719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06231__A1 _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10134_ u_cpu.rf_ram.memory\[32\]\[1\] _04811_ _04815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06042__I _01658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10065_ _04601_ _04456_ _04754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11514__CLK net320 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09859__I0 u_arbiter.i_wb_cpu_rdt\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11664__CLK net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10967_ u_cpu.rf_ram.memory\[85\]\[3\] _05340_ _05342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06137__I2 u_cpu.rf_ram.memory\[118\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06298__A1 _01423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10094__A2 _04572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12706_ u_cpu.cpu.o_wen1 net353 u_cpu.rf_ram_if.wen1_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10898_ _02730_ _05300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10448__B _04602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12637_ _01316_ net63 u_cpu.rf_ram.memory\[24\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12568_ _01247_ net204 u_cpu.rf_ram.memory\[86\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11519_ _00223_ net430 u_cpu.rf_ram.memory\[129\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12499_ _01178_ net37 u_cpu.rf_ram.memory\[107\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout307_I net311 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06661__B _01795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06991_ _01375_ _01371_ _02598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08730_ _03777_ _03779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05942_ u_cpu.cpu.ctrl.o_ibus_adr\[30\] _01560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10403__S _04972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05791__I _01437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08661_ _03733_ _03734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_61_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05873_ u_cpu.cpu.ctrl.o_ibus_adr\[15\] u_cpu.cpu.ctrl.o_ibus_adr\[14\] _01507_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_67_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07722__A1 _01821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07612_ _03000_ _03049_ _03058_ _00161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_93_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08592_ _03676_ _03687_ _03693_ _00506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07543_ _02996_ _03008_ _03015_ _00135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_78_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09475__A1 _04255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07325__I1 u_cpu.rf_ram_if.wdata1_r\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11282__A1 u_cpu.rf_ram.memory\[89\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07474_ _02965_ _02967_ _02968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09213_ _03112_ _04027_ _04090_ _00731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06425_ _01584_ _02040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09144_ _03112_ _02607_ _00709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11034__A1 _05354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09778__A2 _04482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06127__I _01678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06356_ _01619_ _01969_ _01970_ _01971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07789__A1 _02877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10872__I _04829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09075_ u_cpu.rf_ram.memory\[38\]\[5\] _03995_ _03999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06287_ _01735_ _01902_ _01903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08450__A2 _03596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05966__I _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06300__I2 u_cpu.rf_ram.memory\[94\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08026_ u_cpu.rf_ram.memory\[66\]\[6\] _03328_ _03333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08202__A2 _03439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11537__CLK net241 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09950__A2 _04452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09977_ _04626_ _04675_ _00910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08928_ _03902_ _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09173__I _03899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10848__A1 u_cpu.rf_ram.memory\[83\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08859_ _03858_ _03860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06516__A2 _02129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06072__S0 _01686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11870_ _00566_ net516 u_cpu.rf_ram.memory\[136\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10821_ _05209_ _05245_ _05251_ _01178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09466__A1 _04249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08269__A2 _03166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10752_ u_cpu.rf_ram.memory\[79\]\[2\] _05207_ _05208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10683_ _05163_ _05165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09218__A1 u_cpu.rf_ram.memory\[92\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12422_ _01101_ net363 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11025__A1 _03061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09769__A2 _04491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12353_ _01032_ net112 u_cpu.rf_ram.memory\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08441__A2 _03596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11304_ u_cpu.rf_ram.memory\[23\]\[5\] _05551_ _05555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12284_ _00967_ net504 u_arbiter.i_wb_cpu_dbus_adr\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11235_ u_cpu.rf_ram.memory\[98\]\[1\] _05512_ _05514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[60\]_CLK net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12462__CLK net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09941__A2 _04490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11166_ u_cpu.rf_ram.memory\[26\]\[5\] _05469_ _05473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10117_ _04532_ _04710_ _04615_ _04612_ _04801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_11097_ _05425_ _01280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10839__A1 _05206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10048_ _04715_ _04738_ _04740_ _04557_ _00916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_3_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06507__A2 _02120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08628__S _03712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07180__A2 _02753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout257_I net260 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11999_ _00682_ net401 u_cpu.rf_ram.memory\[38\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08427__I _03484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout424_I net434 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11016__A1 _05357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06210_ _01788_ _01827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07190_ _02766_ _02767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06141_ _01739_ _01745_ _01750_ _01756_ _01757_ _01758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_117_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08432__A2 _03590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06072_ u_cpu.rf_ram.memory\[40\]\[0\] u_cpu.rf_ram.memory\[41\]\[0\] u_cpu.rf_ram.memory\[42\]\[0\]
+ u_cpu.rf_ram.memory\[43\]\[0\] _01686_ _01688_ _01689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08162__I _03083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09900_ _04605_ _04606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09917__C1 _04520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[28\]_CLK net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout506 net507 net506 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_8_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09831_ _04451_ _04548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout517 net520 net517 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout528 net530 net528 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XTAP_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout539 net540 net539 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_63_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07943__A1 _03266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09762_ _04475_ _04485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06974_ u_cpu.cpu.alu.i_rs1 _02547_ _02581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05925_ u_cpu.cpu.ctrl.o_ibus_adr\[27\] _01547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08713_ u_cpu.rf_ram.memory\[49\]\[1\] _03767_ _03769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09693_ u_arbiter.i_wb_cpu_rdt\[1\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\]
+ _04417_ _04418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08644_ _03666_ _03722_ _03724_ _00527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05856_ u_arbiter.i_wb_cpu_dbus_adr\[11\] _01493_ _01494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08575_ _03506_ _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05787_ _01435_ u_arbiter.o_wb_cpu_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07526_ _02788_ _03003_ _03004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_74_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09999__A2 _04667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07241__I _02805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08120__A1 _02920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06285__C _01900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06357__S1 _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07457_ _02897_ _02954_ _02957_ _00107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12335__CLK net523 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08671__A2 _03734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09369__S _04186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06408_ _01751_ _02022_ _01755_ _02023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06682__A1 _01876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07388_ _02767_ _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_13_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06109__S1 _01633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09127_ _03111_ _04029_ _04030_ _00704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_06339_ u_cpu.rf_ram.memory\[8\]\[2\] u_cpu.rf_ram.memory\[9\]\[2\] u_cpu.rf_ram.memory\[10\]\[2\]
+ u_cpu.rf_ram.memory\[11\]\[2\] _01574_ _01838_ _01954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06434__A1 _01802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09058_ _03918_ _03988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_123_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08009_ _03270_ _03313_ _03322_ _00294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11020_ _05361_ _05369_ _05376_ _01252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09923__A2 _04627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07934__A1 _03257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06588__I2 u_cpu.rf_ram.memory\[62\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06293__S0 _01747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11922_ _00618_ net153 u_cpu.rf_ram.memory\[12\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07352__S _02879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11853_ _00549_ net510 u_cpu.rf_ram.memory\[137\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09439__A1 _04150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06370__B1 _01982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10804_ _05213_ _05233_ _05240_ _01172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11784_ _00480_ net352 u_cpu.rf_ram.memory\[72\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07151__I _02732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08111__A1 _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10735_ u_cpu.rf_ram.memory\[99\]\[5\] _05192_ _05196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06512__I2 u_cpu.rf_ram.memory\[98\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10666_ _05135_ _05151_ _05154_ _01120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11702__CLK net416 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[50\] u_scanchain_local.module_data_in\[49\] net558 u_arbiter.o_wb_cpu_adr\[12\]
+ net26 u_scanchain_local.module_data_in\[50\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
X_12405_ _01084_ net75 u_cpu.rf_ram.memory\[96\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10218__S _04867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10597_ _03116_ _05111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_86_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12336_ _01016_ net167 u_cpu.rf_ram.memory\[109\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06520__S1 _01908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12267_ _00950_ net521 u_arbiter.i_wb_cpu_dbus_adr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08178__A1 _03412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11218_ _02857_ u_cpu.rf_ram.memory\[0\]\[2\] _05501_ _05504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_9_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12198_ _00881_ net397 u_cpu.rf_ram.memory\[113\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10461__B _04700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11149_ _02777_ _05462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12208__CLK net384 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07326__I _02863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout374_I net375 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09678__A1 _04399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10288__A2 _04907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06690_ _01862_ _02292_ _02301_ _02302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_36_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12358__CLK net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06751__I2 u_cpu.rf_ram.memory\[22\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08360_ _03507_ _03538_ _03546_ _00421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06339__S1 _01838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07311_ _02846_ u_cpu.rf_ram.memory\[1\]\[0\] _02852_ _02853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_60_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08291_ _02766_ _03503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07242_ u_cpu.rf_ram.memory\[81\]\[0\] _02807_ _02808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11382__CLK net185 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06664__A1 _02078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10460__A2 _04520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07173_ _02732_ _02753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06124_ _01673_ _01741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06267__I1 u_cpu.rf_ram.memory\[37\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06967__A2 _02545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06055_ _01671_ _01672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_47_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08169__A1 _02981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09905__A2 _04489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout303 net304 net303 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_119_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout314 net315 net314 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout325 net328 net325 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_86_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06719__A2 _02326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout336 net337 net336 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_119_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09814_ _04504_ _04502_ _04533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout347 net349 net347 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
Xfanout358 net359 net358 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_101_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout369 net372 net369 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_28_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06140__I _01426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09745_ _04446_ _04469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06957_ _02564_ _02565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09669__A1 _04255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05908_ u_cpu.cpu.ctrl.o_ibus_adr\[23\] u_cpu.cpu.ctrl.o_ibus_adr\[22\] _01534_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10279__A2 _04895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09676_ u_arbiter.i_wb_cpu_rdt\[9\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[9\]
+ _01437_ _04401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06888_ _01735_ _02497_ _02498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10597__I _03116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05839_ _01473_ _01478_ _01479_ u_arbiter.o_wb_cpu_adr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08627_ _03714_ _00520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08558_ _03666_ _03668_ _03670_ _00495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07509_ _02903_ _02992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08489_ u_cpu.rf_ram.memory\[140\]\[5\] _03625_ _03629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09841__A1 _01382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06655__A1 _01637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10520_ _05046_ _05060_ _05065_ _01063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10451__A2 _04518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10451_ _04407_ _04518_ _04722_ _05010_ _04469_ _05011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__11875__CLK net519 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10382_ _04827_ _04962_ _04969_ _01021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06958__A2 _01413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12121_ _00804_ net405 u_cpu.rf_ram.memory\[112\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12052_ _00735_ net270 u_cpu.rf_ram.memory\[92\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07907__A1 _03257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11003_ u_cpu.rf_ram.memory\[110\]\[7\] _05348_ _05366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08580__A1 _03684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07383__A2 _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06430__I1 u_cpu.rf_ram.memory\[73\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12500__CLK net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06018__S0 _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08332__A1 _03494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11905_ _00601_ net471 u_cpu.rf_ram.memory\[131\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06894__A1 _02150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11836_ _00532_ net487 u_cpu.rf_ram.memory\[138\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12650__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11767_ _00463_ net479 u_cpu.rf_ram.memory\[140\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08705__I _03509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10718_ _05146_ _05177_ _05185_ _01141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11698_ _00402_ net452 u_cpu.rf_ram.memory\[55\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout122_I net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10649_ u_cpu.rf_ram.memory\[101\]\[4\] _05138_ _05143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09596__B1 _04344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06225__I _01584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09060__A2 _03973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12319_ _00999_ net532 u_cpu.cpu.ctrl.o_ibus_adr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09536__I _03132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08440__I _03497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout491_I net492 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09899__A1 _04549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07860_ _03228_ _03229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_95_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08571__A1 _03678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07374__A2 _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06811_ _01778_ _02421_ _01782_ _02422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_99_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07791_ _03182_ _03184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_42_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12180__CLK net388 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06009__S0 _01622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09530_ _04294_ _04295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06742_ u_cpu.rf_ram.memory\[8\]\[6\] u_cpu.rf_ram.memory\[9\]\[6\] u_cpu.rf_ram.memory\[10\]\[6\]
+ u_cpu.rf_ram.memory\[11\]\[6\] _01591_ _01592_ _02353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10411__S _04983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11748__CLK net256 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08323__A1 _03380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09461_ _03906_ _04247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_58_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06673_ _01697_ _02284_ _02285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10130__A1 u_cpu.rf_ram.memory\[32\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08874__A2 _03860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08412_ _03580_ _00439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09392_ _04204_ _00796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10681__A2 _05162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout35_I u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08343_ _02786_ _03425_ _03536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09823__A1 _04485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11898__CLK net471 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[6\]_CLK net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09823__B2 _04540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06637__A1 _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08274_ _02744_ _03490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07685__I0 _02870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07225_ u_cpu.rf_ram.memory\[21\]\[2\] _02796_ _02797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05860__A2 _01481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07156_ u_cpu.rf_ram_if.wdata0_r\[0\] _02735_ _02737_ _02738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__06135__I _01704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06107_ _01720_ _01722_ _01723_ _01724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07087_ _02673_ _02678_ _01456_ u_arbiter.o_wb_cpu_cyc vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05974__I _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06038_ _01649_ _01654_ _01655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout100 net107 net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_47_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout111 net113 net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_138_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout122 net124 net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_99_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06248__S0 _01863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout133 net139 net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_102_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout144 net145 net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_101_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout155 net156 net155 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout166 net167 net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_25_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06799__S1 _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout177 net184 net177 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_75_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout188 net191 net188 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout199 net201 net199 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_07989_ _03002_ _03310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09728_ _04439_ _04441_ _04453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_60_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08314__A1 _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12673__CLK net289 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09659_ _04244_ _04384_ _04389_ _00878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08865__A2 _03863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06876__A1 _02479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12670_ _01349_ net286 u_cpu.rf_ram.memory\[89\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11621_ _00325_ net101 u_cpu.rf_ram.memory\[29\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08617__A2 _03701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06628__A1 _02147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09130__B _04032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06479__I1 u_cpu.rf_ram.memory\[49\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11552_ _00256_ net253 u_cpu.rf_ram.memory\[76\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10503_ u_cpu.rf_ram.memory\[97\]\[5\] _05047_ _05054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11483_ _00187_ net378 u_cpu.rf_ram_if.rcnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09578__B1 _04331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10434_ _04821_ _04993_ _04999_ _01043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06045__I _01601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10790__I _05231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10365_ _02700_ _02729_ _02847_ _04958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_30_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06800__A1 _01735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12104_ _00787_ net441 u_cpu.rf_ram.memory\[121\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10296_ _04916_ _00988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12035_ _00718_ net313 u_cpu.rf_ram.memory\[91\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06239__S0 _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[13\] u_arbiter.i_wb_cpu_rdt\[10\] net544 u_arbiter.i_wb_cpu_dbus_dat\[7\]
+ net12 u_arbiter.i_wb_cpu_rdt\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_120_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06929__B u_cpu.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10112__A1 _02684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08856__A2 _03848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11126__I _05445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10663__A2 _05152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08636__S _03711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11819_ _00515_ net485 u_cpu.rf_ram.memory\[143\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08608__A2 _03700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout337_I net338 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09281__A2 _04129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06383__C _01711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout504_I net505 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07292__A1 u_cpu.rf_ram.memory\[20\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07010_ u_cpu.cpu.mem_if.signbit _02617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09569__B1 _04321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05842__A2 _01481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11420__CLK net297 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12546__CLK net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05794__I _01440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08961_ _03903_ _03922_ _03927_ _00641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07912_ _03074_ _03262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08892_ _03574_ u_cpu.rf_ram.memory\[12\]\[6\] _03871_ _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08544__A1 _03598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08395__I1 u_cpu.rf_ram.memory\[9\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12696__CLK net379 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07843_ u_cpu.rf_ram.memory\[139\]\[1\] _03217_ _03219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07774_ u_cpu.rf_ram.memory\[40\]\[2\] _03172_ _03173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09513_ _04253_ _04271_ _04279_ _00842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06725_ _01684_ _02336_ _02337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08847__A2 _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09895__I1 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06858__A1 _01772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06656_ u_cpu.rf_ram.memory\[12\]\[5\] u_cpu.rf_ram.memory\[13\]\[5\] u_cpu.rf_ram.memory\[14\]\[5\]
+ u_cpu.rf_ram.memory\[15\]\[5\] _01813_ _01841_ _02268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_80_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09444_ u_cpu.rf_ram.memory\[122\]\[6\] _04230_ _04235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_77_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_75_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10875__I _04832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09375_ _04192_ u_cpu.rf_ram.memory\[8\]\[3\] _04186_ _04193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06587_ _01569_ _02199_ _01867_ _02200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_127_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12076__CLK net318 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08326_ u_cpu.rf_ram.memory\[54\]\[0\] _03526_ _03527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06705__S1 _01908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08257_ u_cpu.rf_ram.memory\[57\]\[3\] _03477_ _03479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07208_ _02720_ _02781_ _02782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_105_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08188_ _03423_ _03428_ _03437_ _00358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09024__A2 _03962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07139_ _01658_ _02720_ _02721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_49_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09176__I _03902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07586__A2 _03036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08783__A1 _03759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10150_ _04826_ _04827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10590__A1 _05051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10081_ _04761_ _04762_ _04447_ _04768_ _04769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_82_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[0\]_D net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06749__B _01795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10893__A2 _05290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10983_ _02745_ _05352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12419__CLK net357 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07360__S _02878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07510__A2 _02990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12653_ _01332_ net66 u_cpu.rf_ram.memory\[98\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05879__I _01451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11604_ _00308_ net243 u_cpu.rf_ram.memory\[65\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12584_ _01263_ net207 u_cpu.rf_ram.memory\[87\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11443__CLK net295 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07274__A1 _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11535_ _00239_ net250 u_cpu.rf_ram.memory\[77\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06321__I0 u_cpu.rf_ram.memory\[76\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05824__A2 _01464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09015__A2 _03959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11466_ _00170_ net301 u_cpu.rf_ram.memory\[50\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10417_ _04196_ u_cpu.rf_ram.memory\[2\]\[5\] _04982_ _04989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10226__S _04867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11397_ _00101_ net299 u_cpu.rf_ram.memory\[42\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07577__A2 _03036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11593__CLK net244 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08774__A1 _03750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06503__I _01665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10348_ u_cpu.cpu.ctrl.o_ibus_adr\[26\] _04943_ _04945_ _01547_ _04947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_98_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10581__A1 _05039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10279_ _04833_ _04895_ _04904_ _00983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.out_flop_D u_scanchain_local.module_data_in\[69\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08526__A1 _03600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12018_ _00701_ net450 u_cpu.rf_ram.memory\[36\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout287_I net288 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06632__S0 _01798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10884__A2 _05289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07334__I _02869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout454_I net455 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08829__A2 _03839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06510_ _02008_ _02123_ _02124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12099__CLK net448 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10636__A2 _05133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07490_ u_cpu.rf_ram.memory\[45\]\[6\] _02973_ _02978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07501__A2 _02984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06441_ u_cpu.rf_ram.memory\[140\]\[2\] u_cpu.rf_ram.memory\[141\]\[2\] u_cpu.rf_ram.memory\[142\]\[2\]
+ u_cpu.rf_ram.memory\[143\]\[2\] _01820_ _01821_ _02056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09160_ _03982_ _04045_ _04052_ _00715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06372_ _01876_ _01986_ _01987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08165__I _03086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09254__A2 _04106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08111_ _03345_ _03382_ _03388_ _00330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09091_ u_cpu.rf_ram.memory\[37\]\[3\] _04007_ _04009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07265__A1 _02746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08042_ _03342_ _03337_ _03344_ _00305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06863__I1 u_cpu.rf_ram.memory\[33\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11936__CLK net462 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09006__A2 _03950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07017__A1 _02612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10947__I0 _04192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07509__I _02903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08765__A1 _03761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09993_ _04688_ _04689_ _04619_ _04690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10572__A1 _04713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06240__A2 _01855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08944_ _02771_ _03915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08517__A1 _03588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08875_ u_cpu.rf_ram.memory\[130\]\[7\] _03858_ _03869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06623__S0 _02142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07826_ u_cpu.rf_ram.memory\[129\]\[2\] _03208_ _03209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07740__A2 _03146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07757_ _03078_ _03154_ _03161_ _00203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10088__B1 _04443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06708_ _01691_ _02319_ _01709_ _02320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07688_ _03110_ _00185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09427_ _03180_ _04224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11466__CLK net301 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06639_ _01791_ _02251_ _01805_ _02252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_9_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09358_ _04154_ _04174_ _04181_ _00785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09245__A2 _04109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07256__A1 _02773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08309_ _03491_ _03513_ _03516_ _00400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09289_ u_cpu.rf_ram.memory\[117\]\[5\] _04133_ _04137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11320_ _03119_ _05563_ _05564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11251_ _05522_ _05523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09953__B1 _04652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10202_ u_arbiter.i_wb_cpu_dbus_adr\[11\] u_arbiter.i_wb_cpu_dbus_adr\[10\] _04855_
+ _04859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11182_ u_cpu.rf_ram.memory\[25\]\[3\] _05481_ _05483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10563__A1 u_cpu.rf_ram.memory\[96\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10133_ _04813_ _04814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06231__A2 _01846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10064_ _04532_ _04709_ _04753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_62_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[6\] u_arbiter.i_wb_cpu_rdt\[3\] net548 u_arbiter.i_wb_cpu_dbus_dat\[0\]
+ net15 u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_75_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12241__CLK net260 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07154__I _02726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09859__I1 u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10966_ _05275_ _05336_ _05341_ _01233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09484__A2 _04262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06137__I3 u_cpu.rf_ram.memory\[119\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12705_ u_cpu.cpu.o_wen0 net353 u_cpu.rf_ram_if.wen0_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06298__A2 _01901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06542__I0 u_cpu.rf_ram.memory\[64\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10897_ _05286_ _05290_ _05299_ _01206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_12636_ _01315_ net63 u_cpu.rf_ram.memory\[24\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_u_scanchain_local.scan_flop\[33\]_D u_arbiter.i_wb_cpu_rdt\[30\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11043__A2 _05379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12567_ _01246_ net163 u_cpu.rf_ram.memory\[110\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10251__B1 _04886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08995__A1 u_cpu.rf_ram.memory\[125\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11518_ _00222_ net321 u_cpu.rf_ram.memory\[119\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10464__B _05022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12498_ _01177_ net38 u_cpu.rf_ram.memory\[107\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout202_I net209 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11449_ _00153_ net299 u_cpu.rf_ram.memory\[43\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08747__A1 _03763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06233__I _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06990_ u_cpu.cpu.state.init_done _02597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11339__CLK net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05941_ _01489_ _01558_ _01559_ u_arbiter.o_wb_cpu_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09172__A1 _04056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05872_ _01502_ _01499_ u_cpu.cpu.ctrl.o_ibus_adr\[15\] _01506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08660_ _02876_ _02940_ _03733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06376__I3 u_cpu.rf_ram.memory\[39\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07611_ u_cpu.rf_ram.memory\[48\]\[7\] _03047_ _03058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08591_ u_cpu.rf_ram.memory\[70\]\[3\] _03691_ _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07542_ u_cpu.rf_ram.memory\[51\]\[5\] _03011_ _03015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09475__A2 _04240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07473_ _02966_ _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_126_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09212_ _02597_ _04038_ _04090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06424_ _01683_ _02039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_u_scanchain_local.scan_flop\[24\]_D u_arbiter.i_wb_cpu_rdt\[21\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09227__A2 _04097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09143_ _04042_ _00708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11034__A2 _05380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06355_ _01602_ _01970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07789__A2 _03181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09074_ _03982_ _03991_ _03998_ _00683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08623__I _03711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06286_ u_cpu.rf_ram.memory\[124\]\[1\] u_cpu.rf_ram.memory\[125\]\[1\] u_cpu.rf_ram.memory\[126\]\[1\]
+ u_cpu.rf_ram.memory\[127\]\[1\] _01736_ _01737_ _01902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_11_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10793__A1 _05199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08025_ _03266_ _03325_ _03332_ _00300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10093__C _04511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08738__A1 u_cpu.rf_ram.memory\[136\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06143__I _01565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10545__A1 u_cpu.rf_ram.memory\[95\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07410__A1 _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09976_ u_cpu.cpu.immdec.imm30_25\[1\] _04672_ _04674_ u_cpu.cpu.immdec.imm30_25\[2\]
+ _04675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_89_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05982__I _01584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09454__I _03899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08927_ _02750_ _03902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05972__A1 _01580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09163__A1 u_cpu.rf_ram.memory\[91\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08858_ _03858_ _03859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07713__A2 _01386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08910__A1 u_cpu.rf_ram.memory\[22\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07809_ _03195_ _03184_ _03196_ _00220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06072__S1 _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08789_ _03201_ _03814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10820_ u_cpu.rf_ram.memory\[107\]\[3\] _05249_ _05251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09466__A2 _04239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10751_ _05200_ _05207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_41_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[15\]_D u_arbiter.i_wb_cpu_rdt\[12\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06318__I _01612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10682_ _05163_ _05164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_13_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12421_ _01100_ net358 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07229__A1 u_cpu.rf_ram.memory\[21\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11025__A2 _05243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12352_ _01031_ net135 u_cpu.rf_ram.memory\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10784__A1 _05213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11303_ _02906_ _05547_ _05554_ _01357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12283_ _00966_ net504 u_arbiter.i_wb_cpu_dbus_adr\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07149__I _02730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12607__CLK net380 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11234_ _05444_ _05511_ _05513_ _01329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11165_ _05456_ _05465_ _05472_ _01301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10116_ _04772_ _04796_ _04799_ _04800_ _00924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_27_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11096_ _05424_ u_cpu.cpu.genblk3.csr.mcause3_0\[1\] _05417_ _05425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_49_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10047_ u_cpu.cpu.immdec.imm19_12_20\[1\] _04636_ _04739_ _04740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_62_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10839__A2 _05257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08901__A1 u_cpu.rf_ram.memory\[22\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11781__CLK net236 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11998_ _00681_ net400 u_cpu.rf_ram.memory\[38\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09701__I0 u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07468__A1 _02913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout152_I net154 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10949_ _04194_ u_cpu.rf_ram.memory\[10\]\[4\] _05326_ _05331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_90_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11264__A2 _05527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11134__I _05445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11016__A2 _05368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12137__CLK net403 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12619_ _01298_ net52 u_cpu.rf_ram.memory\[26\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06691__A2 _02274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06140_ _01426_ _01757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08443__I _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10775__A1 _05204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06071_ _01687_ _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_126_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12287__CLK net502 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09917__C2 _04608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10527__A1 u_cpu.rf_ram.memory\[94\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09830_ _04427_ _04546_ _04491_ _04547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xfanout507 net537 net507 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout518 net519 net518 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XTAP_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout529 net530 net529 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07943__A2 _03275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09761_ _04470_ _04484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06597__I3 u_cpu.rf_ram.memory\[39\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06973_ _02577_ _02580_ u_cpu.cpu.o_wdata1 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09145__A1 _01432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08712_ _03745_ _03766_ _03768_ _00551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05924_ _01524_ _01545_ _01546_ u_arbiter.o_wb_cpu_adr\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09692_ _04413_ _04417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_fanout65_I net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08643_ u_cpu.rf_ram.memory\[138\]\[0\] _03723_ _03724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05855_ _01451_ _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_66_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08574_ _03680_ _03669_ _03681_ _00500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05786_ _01431_ _01434_ _01435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07525_ u_cpu.cpu.immdec.imm11_7\[2\] u_cpu.cpu.immdec.imm11_7\[3\] _02724_ _03003_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07459__A1 u_cpu.rf_ram.memory\[46\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11255__A2 _05524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10088__C _04553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08120__A2 _03005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06138__I _01662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07456_ u_cpu.rf_ram.memory\[46\]\[1\] _02955_ _02957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06407_ u_cpu.rf_ram.memory\[116\]\[2\] u_cpu.rf_ram.memory\[117\]\[2\] u_cpu.rf_ram.memory\[118\]\[2\]
+ u_cpu.rf_ram.memory\[119\]\[2\] _01752_ _01753_ _02022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07387_ _02907_ _02893_ _02908_ _00086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09126_ u_cpu.cpu.state.o_cnt\[2\] _02563_ _04030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_13_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11504__CLK net295 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06338_ _01564_ _01889_ _01953_ _00001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_109_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06434__A2 _02048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06269_ u_cpu.rf_ram.memory\[32\]\[1\] u_cpu.rf_ram.memory\[33\]\[1\] u_cpu.rf_ram.memory\[34\]\[1\]
+ u_cpu.rf_ram.memory\[35\]\[1\] _01705_ _01707_ _01885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09057_ _03986_ _03973_ _03987_ _00677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06985__A3 _01386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08008_ u_cpu.rf_ram.memory\[67\]\[7\] _03311_ _03322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11654__CLK net220 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11191__A1 _05462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07934__A2 _03274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06588__I3 u_cpu.rf_ram.memory\[63\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09959_ _04546_ _04603_ _04659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06293__S1 _01908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09136__A1 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09687__A2 _04411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11921_ _00617_ net150 u_cpu.rf_ram.memory\[12\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07698__A1 _03112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11852_ _00548_ net509 u_cpu.rf_ram.memory\[137\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09439__A2 _04226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06370__A1 _01978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10803_ u_cpu.rf_ram.memory\[106\]\[5\] _05236_ _05240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11246__A2 _05515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11783_ _00479_ net352 u_cpu.rf_ram.memory\[72\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10734_ _05142_ _05188_ _05195_ _01147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06048__I _01397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06122__A1 _01735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06512__I3 u_cpu.rf_ram.memory\[99\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07870__A1 _03191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06673__A2 _02284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10665_ u_cpu.rf_ram.memory\[102\]\[1\] _05152_ _05154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12404_ _01083_ net74 u_cpu.rf_ram.memory\[96\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10596_ _05057_ _05101_ _05110_ _01094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_12335_ _01015_ net523 u_cpu.cpu.ctrl.o_ibus_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xu_scanchain_local.scan_flop\[43\] u_scanchain_local.module_data_in\[42\] net559 u_arbiter.o_wb_cpu_adr\[5\]
+ net27 u_scanchain_local.module_data_in\[43\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12266_ _00949_ net521 u_arbiter.i_wb_cpu_dbus_adr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11217_ _05503_ _01322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06808__S0 _01798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06189__A1 _01802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12197_ _00880_ net396 u_cpu.rf_ram.memory\[113\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10461__C _04581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07925__A2 _03253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06511__I _01673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11148_ _05460_ _05447_ _05461_ _01295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09127__A1 _03111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11079_ u_cpu.rf_ram.memory\[88\]\[5\] _05408_ _05412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09678__A2 _04400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout367_I net394 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06200__I2 u_cpu.rf_ram.memory\[138\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout534_I net535 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07310_ _02851_ _02852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_36_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11527__CLK net488 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08290_ _03501_ _03487_ _03502_ _00395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07241_ _02805_ _02807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10409__S _04983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07172_ _02751_ _02752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10748__A1 u_cpu.rf_ram.memory\[79\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06123_ _01671_ _01740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11677__CLK net286 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06054_ _01567_ _01671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08169__A2 _03425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08413__I0 _03564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout304 net305 net304 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout315 net323 net315 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout326 net328 net326 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
X_09813_ _04411_ _04478_ _04532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_87_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07916__A2 _03260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout337 net338 net337 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_100_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout348 net349 net348 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_28_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout359 net366 net359 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__09118__A1 _03986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09744_ _04425_ _04468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06956_ u_cpu.cpu.mem_bytecnt\[1\] u_cpu.cpu.state.o_cnt\[2\] u_cpu.cpu.mem_bytecnt\[0\]
+ _02564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_28_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09732__I _04456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09669__A2 _04385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05907_ u_cpu.cpu.ctrl.o_ibus_adr\[23\] _01531_ _01533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_41_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09675_ u_arbiter.i_wb_cpu_rdt\[10\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[10\]
+ _01438_ _04400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_36_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06887_ u_cpu.rf_ram.memory\[92\]\[7\] u_cpu.rf_ram.memory\[93\]\[7\] u_cpu.rf_ram.memory\[94\]\[7\]
+ u_cpu.rf_ram.memory\[95\]\[7\] _02142_ _01688_ _02497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08626_ _03564_ u_cpu.rf_ram.memory\[14\]\[1\] _03712_ _03714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05838_ u_arbiter.i_wb_cpu_dbus_adr\[8\] _01461_ _01479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06352__A1 _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10099__B _04550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08557_ u_cpu.rf_ram.memory\[71\]\[0\] _03669_ _03670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05769_ u_cpu.cpu.immdec.imm19_12_20\[7\] _01367_ _01420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07508_ _02989_ _02984_ _02991_ _00124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08488_ _03600_ _03621_ _03628_ _00467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09841__A2 _04396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06655__A2 _02266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07439_ u_cpu.rf_ram.memory\[42\]\[2\] _02946_ _02947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10450_ _04763_ _05009_ _04560_ _05010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_109_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09109_ u_cpu.rf_ram.memory\[36\]\[2\] _04019_ _04020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07604__A1 _02992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10381_ u_cpu.rf_ram.memory\[109\]\[5\] _04965_ _04969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12120_ _00803_ net137 u_cpu.rf_ram.memory\[11\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08811__I _03506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09357__A1 u_cpu.rf_ram.memory\[121\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08404__I0 _03574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12051_ _00734_ net270 u_cpu.rf_ram.memory\[92\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09843__S _01447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[52\]_SE net561 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07907__A2 _03254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11002_ _02777_ _05365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06331__I _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05918__A1 u_cpu.cpu.ctrl.o_ibus_adr\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09109__A1 u_cpu.rf_ram.memory\[36\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06591__A1 _02098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06018__S1 _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08332__A2 _03525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11904_ _00600_ net458 u_cpu.rf_ram.memory\[131\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06733__I3 u_cpu.rf_ram.memory\[143\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11835_ _00531_ net485 u_cpu.rf_ram.memory\[138\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[27\]_CLK net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08096__A1 _03351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11766_ _00462_ net512 u_cpu.rf_ram.memory\[141\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10978__A1 _02920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10717_ u_cpu.rf_ram.memory\[104\]\[6\] _05180_ _05185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06646__A2 _02258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11697_ _00401_ net452 u_cpu.rf_ram.memory\[55\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07111__B _02696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10648_ _04823_ _05142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09596__A1 u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout115_I net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10579_ _05099_ _05101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_5_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12318_ _00998_ net529 u_cpu.cpu.ctrl.o_ibus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12249_ _00932_ net272 u_cpu.rf_ram.memory\[32\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11155__A1 u_cpu.rf_ram.memory\[26\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06241__I _01596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout484_I net494 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10902__A1 u_cpu.rf_ram.memory\[84\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06810_ u_cpu.rf_ram.memory\[68\]\[6\] u_cpu.rf_ram.memory\[69\]\[6\] u_cpu.rf_ram.memory\[70\]\[6\]
+ u_cpu.rf_ram.memory\[71\]\[6\] _01779_ _01780_ _02421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_111_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07790_ _03182_ _03183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_95_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06009__S1 _01625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06741_ _01406_ _02303_ _02352_ _00005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_64_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06397__B _01731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08323__A2 _03287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09460_ _04244_ _04239_ _04246_ _00822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08168__I _03004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06672_ u_cpu.rf_ram.memory\[52\]\[5\] u_cpu.rf_ram.memory\[53\]\[5\] u_cpu.rf_ram.memory\[54\]\[5\]
+ u_cpu.rf_ram.memory\[55\]\[5\] _01863_ _01748_ _02284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_91_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12475__CLK net232 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10130__A2 _04811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08411_ _03560_ u_cpu.rf_ram.memory\[15\]\[0\] _03579_ _03580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09391_ _04184_ u_cpu.rf_ram.memory\[11\]\[0\] _04203_ _04204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08342_ _03510_ _03526_ _03535_ _00414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout28_I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08273_ _03485_ _03487_ _03489_ _00391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07834__A1 u_cpu.rf_ram.memory\[129\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08882__I0 _03564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07224_ _02791_ _02796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06416__I _01678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08634__I0 _03572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07155_ u_cpu.rf_ram_if.wdata1_r\[0\] _02736_ _02737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_69_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06106_ _01417_ _01723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07086_ _02597_ _02674_ _02677_ _02678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07062__A2 _02660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06496__S1 _02109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09339__A1 u_cpu.rf_ram.memory\[118\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06037_ u_cpu.rf_ram.memory\[52\]\[0\] u_cpu.rf_ram.memory\[53\]\[0\] u_cpu.rf_ram.memory\[54\]\[0\]
+ u_cpu.rf_ram.memory\[55\]\[0\] _01651_ _01653_ _01654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_102_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout101 net104 net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout112 net113 net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_114_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout123 net124 net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__06151__I _01675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout134 net139 net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__06248__S1 _01653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout145 net147 net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_134_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout156 net157 net156 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout167 net172 net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10602__S _05111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06412__I2 u_cpu.rf_ram.memory\[94\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout178 net180 net178 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_07988_ _03270_ _03300_ _03309_ _00286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06573__A1 _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05990__I _01606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout189 net191 net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09727_ _04451_ _04452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06939_ _02533_ _02547_ _02548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_41_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09511__A1 _04251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08314__A2 _03513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09658_ u_cpu.rf_ram.memory\[113\]\[2\] _04388_ _04389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08078__I _02789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06325__A1 _01914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08609_ _03699_ _03704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09589_ _04341_ _04342_ _00855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11842__CLK net432 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11620_ _00324_ net101 u_cpu.rf_ram.memory\[29\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09814__A2 _04502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11551_ _00255_ net250 u_cpu.rf_ram.memory\[76\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06628__A2 _02240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06479__I2 u_cpu.rf_ram.memory\[50\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10502_ _04826_ _05053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06326__I _01815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11992__CLK net259 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11482_ _00186_ net379 u_cpu.rf_ram_if.rreq_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09578__A1 u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09578__B2 u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10433_ u_cpu.rf_ram.memory\[93\]\[3\] _04997_ _04999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07358__S _02878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07053__A2 _02654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10364_ _04957_ _01015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_87_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12103_ _00786_ net443 u_cpu.rf_ram.memory\[121\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06800__A2 _02410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10295_ u_cpu.cpu.ctrl.o_ibus_adr\[4\] _04915_ _04910_ _01463_ _04916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_78_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07157__I _02738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12034_ _00717_ net319 u_cpu.rf_ram.memory\[91\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06061__I _01417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06239__S1 _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11372__CLK net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09502__A1 _04242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10112__A2 u_cpu.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06867__A2 _02448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08069__A1 _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11818_ _00514_ net485 u_cpu.rf_ram.memory\[143\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07816__A1 _02724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11749_ _00006_ net256 u_cpu.rf_ram.rdata\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout232_I net235 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06236__I _01621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07292__A2 _02837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09569__A1 u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09569__B2 u_arbiter.i_wb_cpu_dbus_dat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08960_ u_cpu.rf_ram.memory\[127\]\[2\] _03926_ _03927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11128__A1 u_cpu.rf_ram.memory\[27\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07911_ _03259_ _03254_ _03261_ _00257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08891_ _03878_ _00620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08544__A2 _03655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07842_ _03179_ _03216_ _03218_ _00231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07773_ _03167_ _03172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11865__CLK net519 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09512_ u_cpu.rf_ram.memory\[33\]\[6\] _04274_ _04279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06724_ u_cpu.rf_ram.memory\[72\]\[5\] u_cpu.rf_ram.memory\[73\]\[5\] u_cpu.rf_ram.memory\[74\]\[5\]
+ u_cpu.rf_ram.memory\[75\]\[5\] _01934_ _01763_ _02336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_65_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10103__A2 _04395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11300__A1 u_cpu.rf_ram.memory\[23\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09443_ _04154_ _04227_ _04234_ _00817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06655_ _01637_ _02266_ _02267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06855__B _01695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09374_ _02860_ _04192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_36_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06586_ u_cpu.rf_ram.memory\[48\]\[4\] u_cpu.rf_ram.memory\[49\]\[4\] u_cpu.rf_ram.memory\[50\]\[4\]
+ u_cpu.rf_ram.memory\[51\]\[4\] _01812_ _02092_ _02199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_36_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07530__I _03006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06574__C _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08325_ _03524_ _03526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_123_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06146__I _01687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08256_ _03412_ _03473_ _03478_ _00385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07207_ u_cpu.raddr\[1\] _02780_ _02781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_14_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08187_ u_cpu.rf_ram.memory\[60\]\[7\] _03426_ _03437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06881__I2 u_cpu.rf_ram.memory\[114\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09457__I _03902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05985__I _01601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07035__A2 _02624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07138_ _02719_ _02720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_88_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09980__A1 _04545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08783__A2 _03803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07069_ u_cpu.rf_ram_if.rdata0\[3\] _02665_ _02666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06794__A1 _01703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11395__CLK net295 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09393__S _04203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10080_ _04763_ _04766_ _04767_ _04658_ _04768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_43_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12640__CLK net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09192__I _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10982_ _05347_ _05349_ _05351_ _01239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06849__A2 _02458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12652_ _01331_ net66 u_cpu.rf_ram.memory\[98\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12020__CLK net379 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09799__A1 _04475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11603_ _00307_ net243 u_cpu.rf_ram.memory\[65\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12583_ _01262_ net169 u_cpu.rf_ram.memory\[111\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11534_ _00238_ net488 u_cpu.rf_ram.memory\[139\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06056__I _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07274__A2 _02819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12170__CLK net383 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11465_ _00169_ net226 u_cpu.rf_ram.memory\[47\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11738__CLK net152 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07026__A2 _02629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10416_ _04988_ _01036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11396_ _00100_ net302 u_cpu.rf_ram.memory\[42\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10030__A1 _04721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09971__A1 u_cpu.cpu.immdec.imm30_25\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08774__A2 _03802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10347_ _04946_ _01009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10306__I _04905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06785__A1 _02008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10278_ u_cpu.rf_ram.memory\[30\]\[7\] _04893_ _04904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09723__A1 _04436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08526__A2 _03643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12017_ _00700_ net450 u_cpu.rf_ram.memory\[36\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_u_scanchain_local.scan_flop\[5\]_CLK net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06632__S1 _02040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout182_I net183 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11137__I _02757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07337__I0 u_cpu.rf_ram_if.wdata1_r\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout447_I net448 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06396__S0 _01729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06440_ _01400_ _02054_ _02055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08446__I _03503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06371_ u_cpu.rf_ram.memory\[40\]\[2\] u_cpu.rf_ram.memory\[41\]\[2\] u_cpu.rf_ram.memory\[42\]\[2\]
+ u_cpu.rf_ram.memory\[43\]\[2\] _01686_ _01688_ _01986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_128_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12513__CLK net203 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08110_ u_cpu.rf_ram.memory\[63\]\[3\] _03386_ _03388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09090_ _03977_ _04003_ _04008_ _00689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07265__A2 _02818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08041_ u_cpu.rf_ram.memory\[65\]\[2\] _03343_ _03344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10417__S _04982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10021__A1 _02675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09962__A1 _04545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08765__A2 _03791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09992_ _04401_ _04452_ _04523_ _04528_ _04617_ _04689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_88_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout95_I net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08943_ _03913_ _03897_ _03914_ _00636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_48_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08517__A2 _03643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05754__B _01401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08874_ _03830_ _03860_ _03868_ _00613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10324__A2 _04929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09190__A2 _04064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07825_ _03203_ _03208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06623__S1 _01915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07756_ u_cpu.rf_ram.memory\[17\]\[4\] _03158_ _03161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05751__A2 _01401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10088__A1 _04401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06707_ u_cpu.rf_ram.memory\[116\]\[5\] u_cpu.rf_ram.memory\[117\]\[5\] u_cpu.rf_ram.memory\[118\]\[5\]
+ u_cpu.rf_ram.memory\[119\]\[5\] _02136_ _01707_ _02319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_71_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07687_ _02873_ u_cpu.rf_ram.memory\[4\]\[7\] _03101_ _03110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06387__S0 _02001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06000__I0 u_cpu.rf_ram.memory\[20\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09426_ _04158_ _04214_ _04223_ _00811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06638_ u_cpu.rf_ram.memory\[76\]\[4\] u_cpu.rf_ram.memory\[77\]\[4\] u_cpu.rf_ram.memory\[78\]\[4\]
+ u_cpu.rf_ram.memory\[79\]\[4\] _02047_ _01793_ _02251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_125_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06700__A1 _02305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07260__I _02817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12193__CLK net403 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09357_ u_cpu.rf_ram.memory\[121\]\[5\] _04177_ _04181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06569_ _01399_ _02181_ _02069_ _02182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_139_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08308_ u_cpu.rf_ram.memory\[55\]\[1\] _03514_ _03516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07256__A2 _02807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09288_ _04068_ _04129_ _04136_ _00760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10260__A1 _03367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08239_ u_cpu.rf_ram.memory\[58\]\[4\] _03465_ _03468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07008__A2 _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11250_ _02830_ _04958_ _05522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08205__A1 u_cpu.rf_ram.memory\[19\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10012__A1 _04505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10201_ _04858_ _00951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09953__A1 _04650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08756__A2 _03794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10126__I _04807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09953__B2 _04653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06606__I2 u_cpu.rf_ram.memory\[106\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11181_ _05451_ _05477_ _05482_ _01307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06767__A1 _02098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06311__S0 _01787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10563__A2 _05088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10132_ _02744_ _04813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10063_ _04553_ _04609_ _04752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_7_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09181__A2 _04064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06909__I3 u_cpu.rf_ram.memory\[143\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07319__I0 _02858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10079__A1 _04407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10796__I _05231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10965_ u_cpu.rf_ram.memory\[85\]\[2\] _05340_ _05341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11410__CLK net224 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12704_ u_cpu.cpu.o_wdata1 net239 u_cpu.rf_ram_if.wdata1_r\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08692__A1 _03752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07495__A2 _02919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06298__A3 _01913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10896_ u_cpu.rf_ram.memory\[69\]\[7\] _05288_ _05299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12635_ _01314_ net63 u_cpu.rf_ram.memory\[24\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10626__I0 u_arbiter.i_wb_cpu_rdt\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11560__CLK net258 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12566_ _01245_ net162 u_cpu.rf_ram.memory\[110\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07247__A2 _02810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12686__CLK net232 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08995__A2 _03947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11517_ _00221_ net400 u_cpu.rf_ram.memory\[119\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10251__B2 _02691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12497_ _01176_ net40 u_cpu.rf_ram.memory\[107\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11448_ _00152_ net299 u_cpu.rf_ram.memory\[43\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09944__A1 _04582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11379_ _00083_ net215 u_cpu.rf_ram.memory\[80\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06302__S0 _01767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06758__A1 _01619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout397_I net399 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05940_ u_arbiter.i_wb_cpu_dbus_adr\[30\] _01493_ _01559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12066__CLK net282 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07345__I _02878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09172__A2 _04058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout564_I net565 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05871_ _01452_ _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07610_ _02998_ _03049_ _03057_ _00160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_93_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08590_ _03673_ _03687_ _03692_ _00505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09560__I _04294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07541_ _02994_ _03007_ _03014_ _00134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07472_ _02782_ _02919_ _02966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_39_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07486__A2 _02973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11903__CLK net457 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09211_ _04089_ _00730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06423_ _02028_ _02032_ _02035_ _02037_ _01925_ _02038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_61_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout10_I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10617__I0 u_arbiter.i_wb_cpu_rdt\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09142_ _04032_ u_cpu.cpu.state.o_cnt_r\[0\] _04042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_33_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08435__A1 _03593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06354_ u_cpu.rf_ram.memory\[16\]\[2\] u_cpu.rf_ram.memory\[17\]\[2\] u_cpu.rf_ram.memory\[18\]\[2\]
+ u_cpu.rf_ram.memory\[19\]\[2\] _01852_ _01968_ _01969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09632__B1 _04295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08986__A2 _03938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09073_ u_cpu.rf_ram.memory\[38\]\[4\] _03995_ _03998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06285_ _01891_ _01894_ _01897_ _01899_ _01900_ _01901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__06997__A1 _02559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10793__A2 _05232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09936__S _01441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08024_ u_cpu.rf_ram.memory\[66\]\[5\] _03328_ _03332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06424__I _01683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08738__A2 _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09935__B2 _04586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06749__A1 _01786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10545__A2 _05076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12409__CLK net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09975_ _04397_ _04666_ _04674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07410__A2 _02925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08926_ _03900_ _03896_ _03901_ _00632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05972__A2 _01586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09163__A2 _04049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08857_ _02722_ _03814_ _03858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12559__CLK net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11433__CLK net326 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07713__A3 _02674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07808_ u_cpu.rf_ram.memory\[119\]\[5\] _03189_ _03196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08910__A2 _03886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08788_ _03484_ _03813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09470__I _03915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[3\]_SE net547 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07739_ _03081_ _03143_ _03150_ _00196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10750_ _04816_ _05206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07477__A2 _02970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08674__A1 u_cpu.rf_ram.memory\[39\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09409_ _04212_ _04214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10681_ _02876_ _05162_ _05163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06780__S0 _02001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12420_ _01099_ net264 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07229__A2 _02796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08814__I _03509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12351_ _01030_ net138 u_cpu.rf_ram.memory\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08977__A2 _03935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06988__A1 _01411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10784__A2 _05221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11302_ u_cpu.rf_ram.memory\[23\]\[4\] _05551_ _05554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12282_ _00965_ net525 u_arbiter.i_wb_cpu_dbus_adr\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11233_ u_cpu.rf_ram.memory\[98\]\[0\] _05512_ _05513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12089__CLK net401 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10536__A2 _05073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11164_ u_cpu.rf_ram.memory\[26\]\[4\] _05469_ _05472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10115_ u_cpu.cpu.immdec.imm19_12_20\[8\] _04739_ _04800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11095_ _05419_ _05423_ _05424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07165__I _02745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10046_ _04737_ _04739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06599__S0 _01705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08901__A2 _03883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09380__I _02866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06912__A1 _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11997_ _00680_ net400 u_cpu.rf_ram.memory\[38\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07012__S1 u_cpu.cpu.bufreg.lsb\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10948_ _05330_ _01226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08665__A1 u_cpu.rf_ram.memory\[39\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06515__I1 u_cpu.rf_ram.memory\[125\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10472__A1 _04525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout145_I net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10879_ _05288_ _05289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06771__S0 _01721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12618_ _01297_ net52 u_cpu.rf_ram.memory\[26\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09614__B1 _04359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06691__A3 _02283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08968__A2 _03926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12549_ _01228_ net127 u_cpu.rf_ram.memory\[10\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout312_I net315 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09090__A1 _03977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06523__S0 _02136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10775__A2 _05220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06070_ _01623_ _01687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09983__C _04486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09917__A1 _04485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09917__B2 _04599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10527__A2 _05064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout508 net509 net508 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XTAP_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout519 net520 net519 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11456__CLK net370 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09760_ _04467_ _04480_ _04483_ _00885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06972_ _01431_ _02579_ _02580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08711_ u_cpu.rf_ram.memory\[49\]\[0\] _03767_ _03768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05923_ u_arbiter.i_wb_cpu_dbus_adr\[26\] _01539_ _01546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09691_ _04415_ _04416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08642_ _03721_ _03723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05854_ _01485_ _01474_ _01475_ _01491_ _01492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_27_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout58_I net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06847__C _01784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08573_ u_cpu.rf_ram.memory\[71\]\[5\] _03674_ _03681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05785_ _01433_ _01434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_63_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07524_ _02716_ _02875_ _03002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__07024__B _02629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09853__B1 _04568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10463__A1 _04494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07455_ _02889_ _02954_ _02956_ _00106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06762__S0 _01812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06406_ _01746_ _02020_ _02021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09605__B1 _04344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07386_ u_cpu.rf_ram.memory\[80\]\[4\] _02901_ _02908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09125_ u_cpu.cpu.state.o_cnt\[2\] _02563_ _04029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06337_ _01941_ _01952_ _01953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09081__A1 _02785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12231__CLK net383 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09056_ u_cpu.rf_ram.memory\[123\]\[6\] _03978_ _03987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06268_ _01882_ _01883_ _01884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09908__A1 _04399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08007_ _03268_ _03313_ _03321_ _00293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06199_ _01815_ _01816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05993__I _01609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07395__A1 _02913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12381__CLK net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11191__A2 _05478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09958_ _04470_ _04485_ _04658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11949__CLK net461 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09136__A2 _04026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08909_ _03826_ _03882_ _03889_ _00627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07147__A1 u_cpu.cpu.immdec.imm11_7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09889_ u_cpu.rf_ram.memory\[114\]\[6\] _04592_ _04597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11920_ _00616_ net150 u_cpu.rf_ram.memory\[12\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07698__A2 _03119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11851_ _00547_ net508 u_cpu.rf_ram.memory\[137\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06370__A2 _01980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10802_ _05211_ _05232_ _05239_ _01171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11782_ _00478_ net237 u_cpu.rf_ram.memory\[13\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09695__I0 u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10454__A1 _04398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10733_ u_cpu.rf_ram.memory\[99\]\[4\] _05192_ _05195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06122__A2 _01738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06753__S0 _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11329__CLK net217 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10664_ _05130_ _05151_ _05153_ _01119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07870__A2 _03229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12403_ _01082_ net74 u_cpu.rf_ram.memory\[96\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05881__A1 _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09072__A1 _03980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10595_ u_cpu.rf_ram.memory\[28\]\[7\] _05099_ _05110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12334_ _01014_ net523 u_cpu.cpu.ctrl.o_ibus_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06064__I _01426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11479__CLK net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06681__I0 u_cpu.rf_ram.memory\[40\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[36\] u_scanchain_local.module_data_in\[35\] net556 u_arbiter.i_wb_cpu_dbus_dat\[30\]
+ net24 u_scanchain_local.module_data_in\[36\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
X_12265_ _00948_ net515 u_arbiter.i_wb_cpu_dbus_adr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10509__A2 _05040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11216_ _02854_ u_cpu.rf_ram.memory\[0\]\[1\] _05501_ _05503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_64_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06808__S1 _02040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12196_ _00879_ net396 u_cpu.rf_ram.memory\[113\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07386__A1 u_cpu.rf_ram.memory\[80\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11182__A2 _05481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11147_ u_cpu.rf_ram.memory\[27\]\[6\] _05452_ _05461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05936__A2 _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11078_ _05359_ _05404_ _05411_ _01275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09678__A3 _04401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10029_ _04409_ _04549_ _04434_ _04723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_36_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07623__I _03067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout262_I net266 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12104__CLK net441 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout527_I net535 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06744__S0 _01813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07240_ _02805_ _02806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12254__CLK net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07171_ _02750_ _02751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06122_ _01735_ _01738_ _01739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08810__A1 _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06267__I3 u_cpu.rf_ram.memory\[39\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06053_ _01666_ _01669_ _01670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout305 net306 net305 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout316 net317 net316 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_87_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09812_ _02557_ _04396_ _04531_ _00889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout327 net328 net327 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_141_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout338 net395 net338 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout349 net355 net349 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_113_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09743_ _04466_ _04467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06955_ u_cpu.cpu.state.o_cnt_r\[3\] _02563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07129__A1 _02708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05906_ _01505_ _01530_ _01531_ _01532_ u_arbiter.o_wb_cpu_adr\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_100_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09674_ u_arbiter.i_wb_cpu_rdt\[11\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[11\]
+ _01437_ _04399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06886_ _01647_ _02486_ _02495_ _02496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_55_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08625_ _03713_ _00519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05837_ _01476_ _01477_ _01478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06352__A2 _01966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08556_ _03667_ _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06149__I _01671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09677__I0 u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05768_ _01418_ _01419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10436__A1 _04824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07507_ u_cpu.rf_ram.memory\[44\]\[2\] _02990_ _02991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08487_ u_cpu.rf_ram.memory\[140\]\[4\] _03625_ _03628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07301__A1 _02778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06735__S0 _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07438_ _02941_ _02946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08364__I _03548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07852__A2 _03220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09054__A1 _03984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11621__CLK net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07369_ u_cpu.rf_ram.memory\[80\]\[0\] _02894_ _02895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09108_ _04014_ _04019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_109_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08801__A1 _03821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10380_ _04824_ _04961_ _04968_ _01020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07604__A2 _03048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09039_ _03899_ _03975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06663__I0 u_cpu.rf_ram.memory\[20\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11771__CLK net491 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09357__A2 _04177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12050_ _00733_ net270 u_cpu.rf_ram.memory\[92\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06415__I0 u_cpu.rf_ram.memory\[88\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11001_ _05363_ _05350_ _05364_ _01245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11164__A2 _05469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09109__A2 _04019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12127__CLK net407 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08868__A1 _03824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10675__A1 _05144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11903_ _00599_ net457 u_cpu.rf_ram.memory\[131\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12277__CLK net533 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11834_ _00530_ net485 u_cpu.rf_ram.memory\[138\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06059__I _01675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09817__B1 _04525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10427__A1 _04808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11765_ _00461_ net514 u_cpu.rf_ram.memory\[141\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09293__A1 u_cpu.rf_ram.memory\[117\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08096__A2 _03370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06726__S0 _02047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10978__A2 _05243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10716_ _05144_ _05177_ _05184_ _01140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08274__I _02744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07843__A2 _03217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11696_ _00400_ net417 u_cpu.rf_ram.memory\[55\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10309__I _04909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10647_ _05140_ _05132_ _05141_ _01114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09045__A1 _03977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09596__A2 _04347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10578_ _05099_ _05100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_12317_ _00997_ net524 u_cpu.cpu.ctrl.o_ibus_adr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout108_I net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09348__A2 _04174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12248_ _00931_ net272 u_cpu.rf_ram.memory\[32\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06522__I _01704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11155__A2 _05466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10202__I1 u_arbiter.i_wb_cpu_dbus_adr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12179_ _00862_ net387 u_arbiter.i_wb_cpu_dbus_dat\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08020__A2 _03328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10363__B1 _04909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10902__A2 _05303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout477_I net484 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06582__A2 _02194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06740_ _02342_ _02351_ _02352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08449__I _03506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10666__A1 _05135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06671_ _02276_ _02278_ _02280_ _02282_ _01784_ _02283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_08410_ _03578_ _03579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_58_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09390_ _04202_ _04203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_17_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08341_ u_cpu.rf_ram.memory\[54\]\[7\] _03524_ _03535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09284__A1 _04063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11644__CLK net188 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11750__D _00007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06717__S0 _01922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10969__A2 _05340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08272_ u_cpu.rf_ram.memory\[56\]\[0\] _03488_ _03489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07834__A2 _03208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11218__I0 _02857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07223_ _02746_ _02792_ _02795_ _00035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09587__A2 _04338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11794__CLK net352 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07154_ _02726_ _02736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_69_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06105_ u_cpu.rf_ram.memory\[104\]\[0\] u_cpu.rf_ram.memory\[105\]\[0\] u_cpu.rf_ram.memory\[106\]\[0\]
+ u_cpu.rf_ram.memory\[107\]\[0\] _01721_ _01624_ _01722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07085_ _02675_ _02676_ _02677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06270__A1 _01703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06432__I _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09339__A2 _04165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06036_ _01652_ _01653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_47_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08398__I0 _03570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout102 net104 net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_102_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout113 net115 net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout124 net130 net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__10354__B1 _04945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout135 net137 net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_47_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09743__I _04466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout146 net147 net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_102_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout157 net158 net157 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout168 net170 net168 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_47_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07987_ u_cpu.rf_ram.memory\[68\]\[7\] _03298_ _03309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout179 net183 net179 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06573__A2 _02185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07770__A1 _03060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09726_ _04439_ _04450_ _04451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06938_ _02546_ _02547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_60_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09511__A2 _04271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09657_ _04383_ _04388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06869_ _02117_ _02478_ _02479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08608_ _03671_ _03700_ _03703_ _00512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09588_ u_arbiter.i_wb_cpu_rdt\[11\] _04334_ _04331_ u_arbiter.i_wb_cpu_dbus_dat\[11\]
+ _04342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08539_ _03593_ _03655_ _03658_ _00488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_19_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09275__A1 _02785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11550_ _00254_ net261 u_cpu.rf_ram.memory\[74\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11082__A1 _05363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10501_ _05051_ _05041_ _05052_ _01057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11481_ _00185_ net133 u_cpu.rf_ram.memory\[4\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10129__I _04809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09027__A1 _03913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09578__A2 _04334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10432_ _04817_ _04993_ _04998_ _01042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06636__I0 u_cpu.rf_ram.memory\[72\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10363_ u_cpu.cpu.ctrl.o_ibus_adr\[31\] _04906_ _04909_ _04956_ _04957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_136_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08250__A2 _03474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12102_ _00785_ net444 u_cpu.rf_ram.memory\[121\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10294_ _04906_ _04915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_111_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08389__I0 _03564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12033_ _00716_ net319 u_cpu.rf_ram.memory\[91\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08002__A2 _03316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11517__CLK net400 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06403__I3 u_cpu.rf_ram.memory\[123\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06564__A2 _02177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07761__A1 _03084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07173__I _02732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11667__CLK net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06867__A3 _02457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07901__I _03253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08069__A2 _03356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11817_ _00513_ net478 u_cpu.rf_ram.memory\[143\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09266__A1 _04066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11073__A1 u_cpu.rf_ram.memory\[88\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11748_ _00005_ net256 u_cpu.rf_ram.rdata\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09018__A1 _03900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout225_I net228 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11679_ _00383_ net314 u_cpu.rf_ram.memory\[57\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07029__B1 _01382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09569__A2 _04326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06680__C _01427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06627__I0 u_cpu.rf_ram.memory\[80\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08241__A2 _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06252__A1 _01656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07910_ u_cpu.rf_ram.memory\[76\]\[2\] _03260_ _03261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08890_ _03572_ u_cpu.rf_ram.memory\[12\]\[5\] _03871_ _03878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10336__B1 _04938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07841_ u_cpu.rf_ram.memory\[139\]\[0\] _03217_ _03218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10887__A1 _05275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12442__CLK net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11745__D _00002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10502__I _04826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07772_ _03068_ _03168_ _03171_ _00208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07083__I _01374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06723_ _01929_ _02334_ _01932_ _02335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09511_ _04251_ _04271_ _04278_ _00841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07504__A1 _02987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09442_ u_cpu.rf_ram.memory\[122\]\[5\] _04230_ _04234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06654_ u_cpu.rf_ram.memory\[8\]\[5\] u_cpu.rf_ram.memory\[9\]\[5\] u_cpu.rf_ram.memory\[10\]\[5\]
+ u_cpu.rf_ram.memory\[11\]\[5\] _01591_ _01838_ _02266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA_fanout40_I net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09373_ _04191_ _00790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06585_ _01697_ _02197_ _02198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11064__A1 _05365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08324_ _03524_ _03525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05818__A1 _01456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09009__A1 _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08255_ u_cpu.rf_ram.memory\[57\]\[2\] _03477_ _03478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08480__A2 _03622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06871__B _01587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07206_ u_cpu.rf_ram_if.rcnt\[1\] _02717_ u_cpu.raddr\[0\] u_cpu.rf_ram_if.rcnt\[2\]
+ _02780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_88_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06491__A1 _01876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08186_ _03421_ _03428_ _03436_ _00357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07137_ u_cpu.raddr\[0\] _02718_ _02719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_101_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07035__A3 _02640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08232__A2 _03462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09674__S _01437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06162__I _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07068_ _01401_ _02665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06794__A2 _02404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06019_ _01630_ _01635_ _01636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10613__S _05117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[26\]_CLK net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09473__I _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10878__A1 _02785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07743__A1 _03087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09709_ _04429_ _04433_ _04434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_28_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10981_ u_cpu.rf_ram.memory\[110\]\[0\] _05350_ _05351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09496__A1 _02803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09248__A1 _04068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12651_ _01330_ net65 u_cpu.rf_ram.memory\[98\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11602_ _00306_ net243 u_cpu.rf_ram.memory\[65\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12582_ _01261_ net171 u_cpu.rf_ram.memory\[111\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10802__A1 _05211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11533_ _00237_ net488 u_cpu.rf_ram.memory\[139\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08471__A2 _03613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06321__I2 u_cpu.rf_ram.memory\[78\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11464_ _00168_ net226 u_cpu.rf_ram.memory\[47\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09956__C1 _04653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10415_ _04194_ u_cpu.rf_ram.memory\[2\]\[4\] _04983_ _04988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07026__A3 _02602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09420__A1 _04152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11395_ _00099_ net295 u_cpu.rf_ram.memory\[42\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07168__I _02726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10346_ u_cpu.cpu.ctrl.o_ibus_adr\[25\] _04943_ _04945_ u_cpu.cpu.ctrl.o_ibus_adr\[26\]
+ _04946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09971__A2 _04516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07982__A1 _03264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06785__A2 _02395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10277_ _04830_ _04895_ _04903_ _00982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09383__I _02869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12016_ _00699_ net439 u_cpu.rf_ram.memory\[36\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09487__A1 _04247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout175_I net176 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07337__I1 u_cpu.cpu.o_wdata0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11294__A1 _02888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[65\]_SE net554 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10478__B _04487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07631__I _02757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06396__S1 _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout342_I net344 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09239__A1 _04056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11153__I _05464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06370_ _01978_ _01980_ _01982_ _01984_ _01681_ _01985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__06247__I _01650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06691__B _02302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09558__I _04318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08040_ _03336_ _03343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08462__I _03608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09411__A1 _04140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10021__A2 _02703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09962__A2 _04563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09991_ _04497_ _04603_ _04606_ _04688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06615__I3 u_cpu.rf_ram.memory\[123\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07973__A1 _03252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06776__A2 _02386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11832__CLK net478 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08942_ u_cpu.rf_ram.memory\[128\]\[5\] _03904_ _03914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout88_I net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08873_ u_cpu.rf_ram.memory\[130\]\[6\] _03863_ _03868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07824_ _03186_ _03204_ _03207_ _00224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07755_ _03075_ _03154_ _03160_ _00202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11285__A1 _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06706_ _01703_ _02317_ _02318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07686_ _03109_ _00184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06387__S1 _01717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06000__I1 u_cpu.rf_ram.memory\[21\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06637_ _01684_ _02249_ _02250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09425_ u_cpu.rf_ram.memory\[112\]\[7\] _04212_ _04223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12338__CLK net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06157__I _01652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06568_ u_cpu.rf_ram.memory\[12\]\[4\] u_cpu.rf_ram.memory\[13\]\[4\] u_cpu.rf_ram.memory\[14\]\[4\]
+ u_cpu.rf_ram.memory\[15\]\[4\] _01583_ _01841_ _02181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09356_ _04152_ _04173_ _04180_ _00784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06839__I0 u_cpu.rf_ram.memory\[20\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08307_ _03485_ _03513_ _03515_ _00399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07697__B _03118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09287_ u_cpu.rf_ram.memory\[117\]\[4\] _04133_ _04136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08453__A2 _03589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09650__A1 _02803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06499_ _01993_ _02112_ _01996_ _02113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05996__I _01612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11362__CLK net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08238_ _03415_ _03461_ _03467_ _00378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10260__A2 _02921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06854__I3 u_cpu.rf_ram.memory\[59\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08169_ _02981_ _03425_ _03426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10200_ u_arbiter.i_wb_cpu_dbus_adr\[10\] u_arbiter.i_wb_cpu_dbus_adr\[9\] _04855_
+ _04858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10012__A2 _04411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09953__A2 _04510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11180_ u_cpu.rf_ram.memory\[25\]\[2\] _05481_ _05482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06311__S1 _01788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10131_ _04808_ _04810_ _04812_ _00927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_79_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10062_ _04747_ _04748_ _04750_ _04751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07192__A2 _02753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09469__A1 _04251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10079__A2 _04518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11276__A1 _02896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10964_ _05335_ _05340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08141__A1 _02966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12703_ u_cpu.rf_ram_if.wdata1_r\[7\] net235 u_cpu.rf_ram_if.wdata1_r\[6\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08692__A2 _03747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10895_ _05284_ _05290_ _05298_ _01205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06067__I _01683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12634_ _01313_ net63 u_cpu.rf_ram.memory\[24\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[66\] u_scanchain_local.module_data_in\[65\] net554 u_arbiter.o_wb_cpu_adr\[28\]
+ net22 u_scanchain_local.module_data_in\[66\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__08444__A2 _03596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12565_ _01244_ net162 u_cpu.rf_ram.memory\[110\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11516_ _00220_ net400 u_cpu.rf_ram.memory\[119\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12496_ _01175_ net41 u_cpu.rf_ram.memory\[107\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06845__I3 u_cpu.rf_ram.memory\[27\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11447_ _00151_ net300 u_cpu.rf_ram.memory\[43\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10003__A2 _04582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09944__A2 _04641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11378_ _00082_ net187 u_cpu.rf_ram.memory\[80\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06758__A2 _02368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06302__S1 _01768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10329_ _04935_ _01002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07626__I _02751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout292_I net294 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07707__A1 u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05870_ _01501_ _01504_ u_arbiter.o_wb_cpu_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07183__A2 u_cpu.rf_ram_if.wdata0_r\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08380__A1 _03507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout557_I net564 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08507__I0 _03572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06930__A2 u_cpu.cpu.decode.opcode\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05733__A3 u_cpu.cpu.decode.op21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07540_ u_cpu.rf_ram.memory\[51\]\[4\] _03011_ _03014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11267__A1 _02912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08457__I _03608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08132__A1 u_cpu.rf_ram.memory\[62\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07471_ _02939_ _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09210_ _04034_ _02628_ _00710_ _04089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_06422_ _01778_ _02036_ _01782_ _02037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_34_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11385__CLK net217 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10490__A2 _05042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12630__CLK net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09141_ _04039_ _04041_ _00707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10617__I1 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06353_ _01624_ _01968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09632__A1 u_arbiter.i_wb_cpu_rdt\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08435__A2 _03590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09072_ _03980_ _03991_ _03997_ _00682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06284_ _01605_ _01900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_15_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08023_ _03264_ _03324_ _03331_ _00299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08199__A1 u_cpu.rf_ram.memory\[19\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09935__A2 _04629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08920__I _03895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09974_ _04664_ _04671_ _04673_ _00909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12010__CLK net425 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09952__S _01446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08925_ u_cpu.rf_ram.memory\[128\]\[1\] _03897_ _03901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08856_ _03832_ _03848_ _03857_ _00606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09751__I _04431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07174__A2 _02753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07807_ _03080_ _03195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_3639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12160__CLK net311 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05999_ _01615_ _01616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08787_ _03763_ _03803_ _03812_ _00582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11258__A1 u_cpu.rf_ram.memory\[100\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07738_ u_cpu.rf_ram.memory\[16\]\[5\] _03146_ _03150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08123__A1 u_cpu.rf_ram.memory\[62\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09871__A1 _04558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07669_ u_cpu.rf_ram.memory\[50\]\[7\] _03089_ _03100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09871__B2 _04585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09399__S _04203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09408_ _04212_ _04213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_125_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10481__A2 _04630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10680_ _04958_ _05162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_125_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06780__S1 _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11878__CLK net510 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09339_ u_cpu.rf_ram.memory\[118\]\[6\] _04165_ _04170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[4\]_CLK net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12350_ _01029_ net135 u_cpu.rf_ram.memory\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11301_ _02903_ _05547_ _05553_ _01356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_12281_ _00964_ net525 u_arbiter.i_wb_cpu_dbus_adr\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10137__I _04816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11232_ _05510_ _05512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_120_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09926__A2 _04630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07937__A1 _03259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11163_ _05454_ _05465_ _05471_ _01300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10114_ _02676_ _02625_ _04798_ _04799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_27_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06350__I _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11094_ _02684_ _02633_ u_cpu.cpu.genblk3.csr.mcause3_0\[2\] _01386_ _05423_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_103_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10045_ _04737_ _04738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08362__A1 _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11249__A1 _05462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11996_ _00679_ net400 u_cpu.rf_ram.memory\[38\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10947_ _04192_ u_cpu.rf_ram.memory\[10\]\[3\] _05326_ _05330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09862__A1 _04563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10878_ _02785_ _03227_ _05288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06771__S1 _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12674__D _00025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12617_ _01296_ net56 u_cpu.rf_ram.memory\[27\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09614__A1 u_arbiter.i_wb_cpu_rdt\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout138_I net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06525__I _01426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12548_ _01227_ net126 u_cpu.rf_ram.memory\[10\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06979__A2 _02565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12479_ _01158_ net242 u_cpu.rf_ram.memory\[79\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12033__CLK net319 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09917__A2 _04601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07928__A1 _03272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout509 net510 net509 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06260__I _01683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06971_ _02578_ _02579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12183__CLK net389 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08710_ _03765_ _03767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05922_ u_cpu.cpu.ctrl.o_ibus_adr\[26\] _01544_ _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09690_ _03114_ u_arbiter.i_wb_cpu_rdt\[0\] _04414_ _04415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_41_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09571__I _04327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05853_ u_cpu.cpu.ctrl.o_ibus_adr\[11\] u_cpu.cpu.ctrl.o_ibus_adr\[10\] _01491_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08641_ _03721_ _03722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10160__A1 _04833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05784_ _01432_ u_cpu.cpu.state.ibus_cyc _01433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08572_ _03503_ _03680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07523_ _03000_ _02985_ _03001_ _00129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08656__A2 _03726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09853__B2 _04419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07454_ u_cpu.rf_ram.memory\[46\]\[0\] _02955_ _02956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06211__S0 _01826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06405_ u_cpu.rf_ram.memory\[112\]\[2\] u_cpu.rf_ram.memory\[113\]\[2\] u_cpu.rf_ram.memory\[114\]\[2\]
+ u_cpu.rf_ram.memory\[115\]\[2\] _01747_ _01908_ _02020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_50_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06762__S1 _02092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07385_ _02906_ _02907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09605__A1 u_arbiter.i_wb_cpu_rdt\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09605__B2 u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09124_ _04028_ _00703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06336_ _01944_ _01946_ _01949_ _01951_ _01835_ _01952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XANTENNA__05890__A2 _01516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06435__I _01606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09081__A2 _02940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09055_ _03915_ _03986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06267_ u_cpu.rf_ram.memory\[36\]\[1\] u_cpu.rf_ram.memory\[37\]\[1\] u_cpu.rf_ram.memory\[38\]\[1\]
+ u_cpu.rf_ram.memory\[39\]\[1\] _01698_ _01699_ _01883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09746__I _04437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08006_ u_cpu.rf_ram.memory\[67\]\[6\] _03316_ _03321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09908__A2 _04527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06198_ _01706_ _01815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07919__A1 u_cpu.rf_ram.memory\[76\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11400__CLK net293 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12526__CLK net339 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08592__A1 _03676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07395__A2 _02894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07266__I _02817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06170__I _01612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09957_ _04651_ _04656_ _04657_ _00908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_63_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08908_ u_cpu.rf_ram.memory\[22\]\[4\] _03886_ _03889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09888_ _04251_ _04589_ _04596_ _00900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07147__A2 _02724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11550__CLK net261 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08839_ _03846_ _03848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10151__A1 u_cpu.rf_ram.memory\[32\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11850_ _00546_ net508 u_cpu.rf_ram.memory\[137\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10801_ u_cpu.rf_ram.memory\[106\]\[4\] _05236_ _05239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11781_ _00477_ net236 u_cpu.rf_ram.memory\[13\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09695__I1 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10454__A2 _05011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10732_ _05140_ _05188_ _05194_ _01146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06753__S1 _01968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10663_ u_cpu.rf_ram.memory\[102\]\[0\] _05152_ _05153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11251__I _05522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12056__CLK net271 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12402_ _01081_ net75 u_cpu.rf_ram.memory\[96\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10594_ _05055_ _05101_ _05109_ _01093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_12_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12333_ _01013_ net503 u_cpu.cpu.ctrl.o_ibus_adr\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12264_ _00947_ net513 u_arbiter.i_wb_cpu_dbus_adr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06681__I1 u_cpu.rf_ram.memory\[41\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11215_ _05502_ _01321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06269__S0 _01705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12195_ _00878_ net398 u_cpu.rf_ram.memory\[113\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xu_scanchain_local.scan_flop\[29\] u_arbiter.i_wb_cpu_rdt\[26\] net545 u_arbiter.i_wb_cpu_dbus_dat\[23\]
+ net13 u_arbiter.i_wb_cpu_rdt\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_64_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07386__A2 _02901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06080__I _01648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11146_ _02772_ _05460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_7_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11077_ u_cpu.rf_ram.memory\[88\]\[4\] _05408_ _05411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09678__A4 _04402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10028_ _04487_ _04491_ _04722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10330__I _04905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07125__B _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06441__S0 _01820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10693__A2 _05168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout255_I net262 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09835__A1 _04416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11979_ _00019_ net265 u_cpu.rf_ram_if.rdata1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08735__I _03777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06744__S1 _01815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_fanout422_I net423 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07170_ _02735_ u_cpu.rf_ram_if.wdata0_r\[2\] _02749_ _02750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__06255__I _01673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06121_ u_cpu.rf_ram.memory\[124\]\[0\] u_cpu.rf_ram.memory\[125\]\[0\] u_cpu.rf_ram.memory\[126\]\[0\]
+ u_cpu.rf_ram.memory\[127\]\[0\] _01736_ _01737_ _01738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07074__A1 _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12549__CLK net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08810__A2 _03817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06052_ u_cpu.rf_ram.memory\[60\]\[0\] u_cpu.rf_ram.memory\[61\]\[0\] u_cpu.rf_ram.memory\[62\]\[0\]
+ u_cpu.rf_ram.memory\[63\]\[0\] _01639_ _01668_ _01669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_12_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11748__D _00005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10505__I _04829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08574__A1 _03680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11573__CLK net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout306 net338 net306 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_09811_ _04516_ _04530_ _04531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12699__CLK net232 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout317 net322 net317 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_140_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout328 net336 net328 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout339 net340 net339 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_119_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10381__A1 u_cpu.rf_ram.memory\[109\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09742_ _04465_ _04466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_fanout70_I net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06954_ u_cpu.cpu.decode.op22 _02562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07129__A2 _02710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05905_ u_arbiter.i_wb_cpu_dbus_adr\[22\] _01512_ _01532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09673_ _04397_ _04398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06885_ _02488_ _02490_ _02492_ _02494_ _02139_ _02495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_39_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08624_ _03560_ u_cpu.rf_ram.memory\[14\]\[0\] _03712_ _03713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06888__A1 _01735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05836_ _01474_ _01475_ _01477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__10684__A2 _05165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08555_ _03667_ _03668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05767_ _01417_ _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09677__I1 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12079__CLK net319 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07506_ _02983_ _02990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10436__A2 _04993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08486_ _03598_ _03621_ _03627_ _00466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06735__S1 _01616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07437_ _02897_ _02942_ _02945_ _00099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09677__S _01438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06165__I _01627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09054__A2 _03973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07368_ _02892_ _02894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_143_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07065__A1 _01430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09107_ _03975_ _04015_ _04018_ _00696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06319_ u_cpu.rf_ram.memory\[72\]\[1\] u_cpu.rf_ram.memory\[73\]\[1\] u_cpu.rf_ram.memory\[74\]\[1\]
+ u_cpu.rf_ram.memory\[75\]\[1\] _01934_ _01799_ _01935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_30_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07299_ _02773_ _02834_ _02842_ _00064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08801__A2 _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09038_ _03969_ _03972_ _03974_ _00671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08565__A1 _03673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11000_ u_cpu.rf_ram.memory\[110\]\[6\] _05355_ _05364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10372__A1 u_cpu.rf_ram.memory\[109\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06768__C _01427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08868__A2 _03859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10150__I _04826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11902_ _00598_ net459 u_cpu.rf_ram.memory\[132\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10675__A2 _05152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07540__A2 _03011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11833_ _00529_ net478 u_cpu.rf_ram.memory\[138\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09817__A1 _04484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09817__B2 _04535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07679__I0 _02861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10427__A2 _04993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11764_ _00460_ net508 u_cpu.rf_ram.memory\[141\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06726__S1 _01793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10715_ u_cpu.rf_ram.memory\[104\]\[5\] _05180_ _05184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11446__CLK net326 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06351__I0 u_cpu.rf_ram.memory\[20\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11695_ _00399_ net331 u_cpu.rf_ram.memory\[55\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06075__I _01620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10646_ u_cpu.rf_ram.memory\[101\]\[3\] _05138_ _05141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10577_ _05098_ _02982_ _05099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09386__I _02872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11596__CLK net251 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12316_ _00996_ net529 u_cpu.cpu.ctrl.o_ibus_adr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12247_ _00930_ net272 u_cpu.rf_ram.memory\[32\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12178_ _00861_ net386 u_arbiter.i_wb_cpu_dbus_dat\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10363__B2 _04956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11129_ _05444_ _05446_ _05448_ _01289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout372_I net375 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06670_ _01857_ _02281_ _01859_ _02282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10666__A2 _05151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12221__CLK net350 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07531__A2 _03008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06590__I0 u_cpu.rf_ram.memory\[56\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08340_ _03507_ _03526_ _03534_ _00413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09284__A2 _04129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06717__S1 _02151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08271_ _03486_ _03488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07295__A1 _02763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12371__CLK net343 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07222_ u_cpu.rf_ram.memory\[21\]\[1\] _02793_ _02795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07153_ _02734_ _02735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_118_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06104_ _01620_ _01721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__07598__A2 _03049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09992__B1 _04523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07084_ _02532_ _02676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06035_ _01623_ _01652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06270__A2 _01885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08547__A1 u_cpu.rf_ram.memory\[73\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout103 net105 net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout114 net115 net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_141_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout125 net129 net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__10354__B2 u_cpu.cpu.ctrl.o_ibus_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout136 net137 net136 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_113_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout147 net148 net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_25_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout158 net269 net158 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_75_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07986_ _03268_ _03300_ _03308_ _00285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout169 net170 net169 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_68_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07770__A2 _03168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09725_ _03113_ u_arbiter.i_wb_cpu_rdt\[13\] _04449_ _04450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_74_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10106__A1 _04650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06937_ _02541_ _02545_ u_arbiter.i_wb_cpu_dbus_we _02546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06405__S0 _01747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09656_ _04242_ _04384_ _04387_ _00877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06868_ u_cpu.rf_ram.memory\[108\]\[7\] u_cpu.rf_ram.memory\[109\]\[7\] u_cpu.rf_ram.memory\[110\]\[7\]
+ u_cpu.rf_ram.memory\[111\]\[7\] _01639_ _01615_ _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_3_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08607_ u_cpu.rf_ram.memory\[143\]\[1\] _03701_ _03703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05819_ u_cpu.cpu.ctrl.o_ibus_adr\[5\] _01463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11469__CLK net302 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09587_ u_arbiter.i_wb_cpu_dbus_dat\[12\] _04338_ _04341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06799_ u_cpu.rf_ram.memory\[92\]\[6\] u_cpu.rf_ram.memory\[93\]\[6\] u_cpu.rf_ram.memory\[94\]\[6\]
+ u_cpu.rf_ram.memory\[95\]\[6\] _02142_ _01688_ _02410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05999__I _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08538_ u_cpu.rf_ram.memory\[73\]\[1\] _03656_ _03658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09275__A2 _03970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07286__A1 _02740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08469_ u_cpu.rf_ram.memory\[141\]\[5\] _03613_ _03617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10290__B1 _04910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10500_ u_cpu.rf_ram.memory\[97\]\[4\] _05047_ _05052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11480_ _00184_ net142 u_cpu.rf_ram.memory\[4\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09027__A2 _03959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10431_ u_cpu.rf_ram.memory\[93\]\[2\] _04997_ _04998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07589__A2 _03040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09983__B1 _04523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06636__I1 u_cpu.rf_ram.memory\[73\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10362_ _04953_ _04954_ _04955_ _04956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_87_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10593__A1 u_cpu.rf_ram.memory\[28\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12101_ _00784_ net443 u_cpu.rf_ram.memory\[121\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10145__I _02761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10293_ _04914_ _00987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_88_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[3\]_D u_arbiter.i_wb_cpu_rdt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08538__A1 u_cpu.rf_ram.memory\[73\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08389__I1 u_cpu.rf_ram.memory\[9\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12032_ _00715_ net312 u_cpu.rf_ram.memory\[91\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06779__B _02389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12244__CLK net274 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07761__A2 _03155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07513__A2 _02990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11816_ _00512_ net477 u_cpu.rf_ram.memory\[143\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11747_ _00004_ net253 u_cpu.rf_ram.rdata\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05827__A2 _01461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10820__A2 _05249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09018__A2 _03958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11678_ _00382_ net299 u_cpu.rf_ram.memory\[58\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout120_I net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10629_ _05128_ _01109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout218_I net219 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08777__A1 _03752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06533__I _01702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06252__A2 _01866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06883__S0 _02136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08529__A1 u_cpu.rf_ram.memory\[72\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07201__A1 _02734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07840_ _03215_ _03217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10887__A2 _05289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07752__A2 _03158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07771_ u_cpu.rf_ram.memory\[40\]\[1\] _03169_ _03171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11611__CLK net238 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09510_ u_cpu.rf_ram.memory\[33\]\[5\] _04274_ _04278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06722_ u_cpu.rf_ram.memory\[68\]\[5\] u_cpu.rf_ram.memory\[69\]\[5\] u_cpu.rf_ram.memory\[70\]\[5\]
+ u_cpu.rf_ram.memory\[71\]\[5\] _01779_ _01930_ _02334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10639__A2 _05133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08701__A1 _03759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07504__A2 _02984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09441_ _04152_ _04226_ _04233_ _00816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06653_ _01564_ _02216_ _02265_ _00004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_92_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout33_I net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09372_ _04190_ u_cpu.rf_ram.memory\[8\]\[2\] _04186_ _04191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_36_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06584_ u_cpu.rf_ram.memory\[52\]\[4\] u_cpu.rf_ram.memory\[53\]\[4\] u_cpu.rf_ram.memory\[54\]\[4\]
+ u_cpu.rf_ram.memory\[55\]\[4\] _01863_ _01748_ _02197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__11761__CLK net481 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08323_ _03380_ _03287_ _03524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07268__A1 _02752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11064__A2 _05393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08923__I _02744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08254_ _03472_ _03477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09009__A2 _03947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07205_ _02741_ _02778_ _02779_ _00033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08185_ u_cpu.rf_ram.memory\[60\]\[6\] _03431_ _03436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08768__A1 _03201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07136_ u_cpu.rf_ram_if.rcnt\[1\] _02717_ u_cpu.rf_ram_if.rcnt\[2\] _02718_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10575__A1 _03112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07067_ _01430_ _02649_ _02664_ _00009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07440__A1 _02900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12267__CLK net521 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06018_ u_cpu.rf_ram.memory\[28\]\[0\] u_cpu.rf_ram.memory\[29\]\[0\] u_cpu.rf_ram.memory\[30\]\[0\]
+ u_cpu.rf_ram.memory\[31\]\[0\] _01631_ _01634_ _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_102_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10878__A2 _03227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07743__A2 _03143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05754__A1 _01378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07969_ _02831_ _02923_ _03298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09708_ _04431_ _04432_ _04433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_99_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10980_ _05348_ _05350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_95_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09496__A2 _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09639_ u_arbiter.i_wb_cpu_dbus_dat\[29\] _04376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_71_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12650_ _01329_ net65 u_cpu.rf_ram.memory\[98\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09248__A2 _04105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11601_ _00305_ net243 u_cpu.rf_ram.memory\[65\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07259__A1 _02723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12581_ _01260_ net168 u_cpu.rf_ram.memory\[111\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11532_ _00236_ net486 u_cpu.rf_ram.memory\[139\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10802__A2 _05232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06857__I1 u_cpu.rf_ram.memory\[41\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06321__I3 u_cpu.rf_ram.memory\[79\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11463_ _00167_ net226 u_cpu.rf_ram.memory\[47\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08759__A1 _03755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10414_ _04987_ _01035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06353__I _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09956__C2 _04558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10566__A1 _05053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11394_ _00098_ net297 u_cpu.rf_ram.memory\[42\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07431__A1 _02938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10345_ _04908_ _04945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07982__A2 _03299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10276_ u_cpu.rf_ram.memory\[30\]\[6\] _04898_ _04903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09184__A1 u_cpu.rf_ram.memory\[90\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[11\] u_arbiter.i_wb_cpu_rdt\[8\] net544 u_arbiter.i_wb_cpu_dbus_dat\[5\]
+ net12 u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
X_12015_ _00698_ net439 u_cpu.rf_ram.memory\[36\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06617__S0 _02133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07184__I _02761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08931__A1 _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07734__A2 _03146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05745__A1 _01394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06793__I0 u_cpu.rf_ram.memory\[112\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09487__A2 _04258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11784__CLK net352 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07912__I _03074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11294__A2 _05547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout168_I net170 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xserv_1_566 io_oeb[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_94_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10478__C _04575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06528__I _01685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09239__A2 _04105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout335_I net336 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08998__A1 _03900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout502_I net505 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07670__A1 _03087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06263__I _01659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10557__A1 _05044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09990_ _03115_ u_arbiter.i_wb_cpu_rdt\[28\] _04686_ _04687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07973__A2 _03299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08941_ _03912_ _03913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09175__A1 _04061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10513__I _05059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06608__S0 _02122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08872_ _03828_ _03860_ _03867_ _00612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08922__A1 _03894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07823_ u_cpu.rf_ram.memory\[129\]\[1\] _03205_ _03207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07754_ u_cpu.rf_ram.memory\[17\]\[3\] _03158_ _03160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06705_ u_cpu.rf_ram.memory\[112\]\[5\] u_cpu.rf_ram.memory\[113\]\[5\] u_cpu.rf_ram.memory\[114\]\[5\]
+ u_cpu.rf_ram.memory\[115\]\[5\] _02133_ _01908_ _02317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_38_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07489__A1 _02910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07685_ _02870_ u_cpu.rf_ram.memory\[4\]\[6\] _03101_ _03109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_52_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09424_ _04156_ _04214_ _04222_ _00810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06636_ u_cpu.rf_ram.memory\[72\]\[4\] u_cpu.rf_ram.memory\[73\]\[4\] u_cpu.rf_ram.memory\[74\]\[4\]
+ u_cpu.rf_ram.memory\[75\]\[4\] _01934_ _01763_ _02249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06000__I2 u_cpu.rf_ram.memory\[22\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[27\]_D u_arbiter.i_wb_cpu_rdt\[24\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11037__A2 _05384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09355_ u_cpu.rf_ram.memory\[121\]\[4\] _04177_ _04180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06567_ _01637_ _02179_ _02180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08989__A1 _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08306_ u_cpu.rf_ram.memory\[55\]\[0\] _03514_ _03515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06839__I1 u_cpu.rf_ram.memory\[21\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11507__CLK net302 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09286_ _04066_ _04129_ _04135_ _00759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06498_ u_cpu.rf_ram.memory\[32\]\[3\] u_cpu.rf_ram.memory\[33\]\[3\] u_cpu.rf_ram.memory\[34\]\[3\]
+ u_cpu.rf_ram.memory\[35\]\[3\] _01705_ _01994_ _02112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09650__A2 _04224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08237_ u_cpu.rf_ram.memory\[58\]\[3\] _03465_ _03467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07661__A1 u_cpu.rf_ram.memory\[50\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08168_ _03004_ _03425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10548__A1 _05055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07119_ _02695_ _02705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_49_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08099_ _03004_ _03380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10130_ u_cpu.rf_ram.memory\[32\]\[0\] _04811_ _04812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09166__A1 _03988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10061_ _04517_ _04642_ _04749_ _04750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__08213__I0 _02855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08913__A1 _03830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05727__A1 u_cpu.cpu.decode.op21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10720__A1 _05148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06775__I0 u_cpu.rf_ram.memory\[32\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09469__A2 _04240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10963_ _05273_ _05336_ _05339_ _01232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12702_ u_cpu.rf_ram_if.wdata1_r\[6\] net233 u_cpu.rf_ram_if.wdata1_r\[5\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08141__A2 _03005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[18\]_D u_arbiter.i_wb_cpu_rdt\[15\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10894_ u_cpu.rf_ram.memory\[69\]\[6\] _05293_ _05298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12633_ _01312_ net54 u_cpu.rf_ram.memory\[25\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06792__B _01679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10087__I0 u_arbiter.i_wb_cpu_rdt\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12564_ _01243_ net161 u_cpu.rf_ram.memory\[110\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11515_ _00219_ net321 u_cpu.rf_ram.memory\[119\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xu_scanchain_local.scan_flop\[59\] u_scanchain_local.module_data_in\[58\] net562 u_arbiter.o_wb_cpu_adr\[21\]
+ net31 u_scanchain_local.module_data_in\[59\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_89_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12495_ _01174_ net41 u_cpu.rf_ram.memory\[106\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07179__I _02757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11446_ _00150_ net326 u_cpu.rf_ram.memory\[43\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06207__A2 _01822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11200__A2 _05493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11377_ _00081_ net133 u_cpu.rf_ram.memory\[7\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10328_ u_cpu.cpu.ctrl.o_ibus_adr\[18\] _04929_ _04931_ u_cpu.cpu.ctrl.o_ibus_adr\[19\]
+ _04935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09157__A1 u_cpu.rf_ram.memory\[91\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10333__I _04908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10259_ _02672_ _04888_ _04892_ _00975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_79_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[32\]_SE net549 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10011__I0 u_arbiter.i_wb_cpu_rdt\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09952__I0 u_arbiter.i_wb_cpu_rdt\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08904__A1 u_cpu.rf_ram.memory\[22\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout285_I net289 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06766__I0 u_cpu.rf_ram.memory\[56\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08380__A2 _03550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05733__A4 _01372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06930__A3 u_cpu.cpu.branch_op vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11267__A2 _05524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout452_I net455 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07470_ _02916_ _02955_ _02964_ _00113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_78_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06421_ u_cpu.rf_ram.memory\[84\]\[2\] u_cpu.rf_ram.memory\[85\]\[2\] u_cpu.rf_ram.memory\[86\]\[2\]
+ u_cpu.rf_ram.memory\[87\]\[2\] _01922_ _01780_ _02036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_37_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07891__A1 u_cpu.rf_ram.memory\[74\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11019__A2 _05372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09140_ u_cpu.rf_ram_if.rgnt _04040_ _02699_ _04032_ _04041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06352_ _01611_ _01966_ _01967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09632__A2 _04326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10778__A1 _05206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11113__B _04032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06283_ _01728_ _01898_ _01731_ _01899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10508__I _04832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09071_ u_cpu.rf_ram.memory\[38\]\[3\] _03995_ _03997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06207__B _01823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08022_ u_cpu.rf_ram.memory\[66\]\[4\] _03328_ _03331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07817__I _03201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09973_ u_cpu.cpu.immdec.imm30_25\[0\] _04672_ _04673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08924_ _03899_ _03900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08855_ u_cpu.rf_ram.memory\[131\]\[7\] _03846_ _03857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12305__CLK net502 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07806_ _03193_ _03183_ _03194_ _00219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08371__A2 _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08786_ u_cpu.rf_ram.memory\[134\]\[7\] _03801_ _03812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05998_ _01575_ _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11258__A2 _05527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07737_ _03078_ _03142_ _03149_ _00195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08123__A2 _03395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07668_ _03084_ _03091_ _03099_ _00176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09871__A2 _04574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09407_ _02890_ _03970_ _04212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06619_ u_cpu.rf_ram.memory\[116\]\[4\] u_cpu.rf_ram.memory\[117\]\[4\] u_cpu.rf_ram.memory\[118\]\[4\]
+ u_cpu.rf_ram.memory\[119\]\[4\] _02136_ _01753_ _02232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_52_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07599_ _02987_ _03048_ _03051_ _00155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_41_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08383__I _02845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09338_ _04154_ _04162_ _04169_ _00777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10769__A1 _03019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05800__I _01446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07634__A1 _03075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06437__A2 _02038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09269_ u_cpu.rf_ram.memory\[34\]\[5\] _04121_ _04125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11300_ u_cpu.rf_ram.memory\[23\]\[3\] _05551_ _05553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12280_ _00963_ net526 u_arbiter.i_wb_cpu_dbus_adr\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11231_ _05510_ _05511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[55\]_SE net561 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07937__A2 _03274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11162_ u_cpu.rf_ram.memory\[26\]\[3\] _05469_ _05471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10113_ _04511_ _04797_ _04798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10153__I _02771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11093_ _02568_ _05418_ _05422_ _01279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_49_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10044_ _02529_ _04736_ _03117_ _04737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_114_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[4\] u_arbiter.i_wb_cpu_rdt\[1\] net548 u_arbiter.i_wb_cpu_dbus_sel\[2\]
+ net15 u_arbiter.i_wb_cpu_rdt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_76_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06787__B _01663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08362__A2 _03538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11249__A2 _05512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11995_ _00014_ net257 u_cpu.rf_ram_if.rdata0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08114__A2 _03386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06078__I _01678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10946_ _05329_ _01225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09862__A2 _04568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10877_ _05286_ _05271_ _05287_ _01198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11822__CLK net477 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12616_ _01295_ net56 u_cpu.rf_ram.memory\[27\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09614__A2 _04347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12547_ _01226_ net119 u_cpu.rf_ram.memory\[10\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07625__A1 _03068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12478_ _01157_ net190 u_cpu.rf_ram.memory\[79\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12690__D u_cpu.cpu.o_wdata0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08425__I0 _03576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11429_ _00133_ net327 u_cpu.rf_ram.memory\[51\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11185__A1 _05456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07928__A2 _03034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08050__A1 u_cpu.rf_ram.memory\[65\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05939__A1 u_cpu.cpu.ctrl.o_ibus_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10932__A1 _05280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11159__I _05464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12328__CLK net504 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06600__A2 _02212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06970_ _01387_ _02578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_84_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input5_I io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05921_ u_cpu.cpu.ctrl.o_ibus_adr\[25\] _01537_ _01535_ _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08353__A2 _03541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08640_ _02937_ _03698_ _03721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05852_ _01484_ _01486_ u_cpu.cpu.ctrl.o_ibus_adr\[11\] _01490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_54_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11352__CLK net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10160__A2 _04811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07372__I _02896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08571_ _03678_ _03668_ _03679_ _00499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05783_ net2 _01432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_54_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08105__A2 _03383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07522_ u_cpu.rf_ram.memory\[44\]\[7\] _02983_ _03001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09853__A2 _04566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07453_ _02953_ _02955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06211__S1 _01827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06404_ _01904_ _02018_ _01744_ _02019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_37_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07384_ _02762_ _02906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09605__A2 _04347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09123_ _03111_ _04027_ _04028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_109_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06335_ _01830_ _01950_ _01419_ _01951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09054_ _03984_ _03973_ _03985_ _00676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07092__A2 _02616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06266_ _01665_ _01882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08005_ _03266_ _03313_ _03320_ _00292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06197_ _01813_ _01814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_11_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11176__A1 _05444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07919__A2 _03260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10923__A1 _05268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09956_ u_cpu.cpu.immdec.imm24_20\[4\] _04628_ _04633_ u_cpu.cpu.immdec.imm30_25\[0\]
+ _04653_ _04558_ _04657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_28_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09762__I _04475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08907_ _03824_ _03882_ _03888_ _00626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09887_ u_cpu.rf_ram.memory\[114\]\[5\] _04592_ _04596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09541__A1 u_arbiter.i_wb_cpu_dbus_dat\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08838_ _03846_ _03847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08769_ _03801_ _03802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11845__CLK net432 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10800_ _05209_ _05232_ _05238_ _01170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11780_ _00476_ net145 u_cpu.rf_ram.memory\[13\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10731_ u_cpu.rf_ram.memory\[99\]\[3\] _05192_ _05194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07855__A1 _03197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10662_ _05150_ _05152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11995__CLK net257 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05961__S0 _01574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12401_ _01080_ net75 u_cpu.rf_ram.memory\[96\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10593_ u_cpu.rf_ram.memory\[28\]\[6\] _05104_ _05109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12332_ _01012_ net501 u_cpu.cpu.ctrl.o_ibus_adr\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12263_ _00946_ net513 u_arbiter.i_wb_cpu_dbus_adr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08407__I0 _03576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06681__I2 u_cpu.rf_ram.memory\[42\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11167__A1 _05458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11214_ _02845_ u_cpu.rf_ram.memory\[0\]\[0\] _05501_ _05502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06269__S1 _01707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12194_ _00877_ net403 u_cpu.rf_ram.memory\[113\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10914__A1 _05282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11145_ _05458_ _05447_ _05459_ _01294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11375__CLK net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06594__A1 _01876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12620__CLK net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11076_ _05357_ _05404_ _05410_ _01274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08335__A2 _03529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10027_ _04404_ u_arbiter.i_wb_cpu_rdt\[7\] _04720_ _04721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_3_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08288__I _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06346__A1 _01958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06897__A2 _02506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06441__S1 _01821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11978_ _00018_ net265 u_cpu.rf_ram_if.rdata1\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09835__A2 _04472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12685__D u_cpu.rf_ram_if.wdata0_r\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10929_ u_cpu.rf_ram.memory\[59\]\[3\] _05318_ _05320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08894__I0 _03576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout248_I net267 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12000__CLK net401 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06536__I _01609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout415_I net417 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06120_ _01687_ _01737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07074__A2 _02656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06121__I1 u_cpu.rf_ram.memory\[125\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06051_ _01667_ _01668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11158__A1 _05449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11718__CLK net415 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08023__A1 _03264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10905__A1 _05273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10007__B _04619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09810_ _04518_ _04520_ _04524_ _04525_ _04529_ _04530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_87_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout307 net311 net307 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_114_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09771__A1 _03118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout318 net322 net318 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout329 net332 net329 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_98_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10381__A2 _04965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09741_ _04464_ _04465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06953_ _01380_ _01383_ _02561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_39_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09523__A1 _04285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08326__A2 _03526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[3\]_CLK net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05904_ _01528_ _01529_ _01531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09672_ _03117_ _04397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06884_ _01691_ _02493_ _01709_ _02494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_fanout63_I net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08623_ _03711_ _03712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05835_ _01474_ _01475_ _01476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08554_ _02876_ _03227_ _03667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05766_ _01407_ _01416_ _01417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_58_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07505_ _02899_ _02989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07837__A1 _03199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08485_ u_cpu.rf_ram.memory\[140\]\[3\] _03625_ _03627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06446__I _01613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07436_ u_cpu.rf_ram.memory\[42\]\[1\] _02943_ _02945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07367_ _02892_ _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06890__B _01744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09106_ u_cpu.rf_ram.memory\[36\]\[1\] _04016_ _04018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06318_ _01612_ _01934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08262__A1 _03419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07298_ u_cpu.rf_ram.memory\[20\]\[6\] _02837_ _02842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09037_ u_cpu.rf_ram.memory\[123\]\[0\] _03973_ _03974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06249_ _01649_ _01864_ _01865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06663__I2 u_cpu.rf_ram.memory\[22\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11398__CLK net301 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09693__S _04417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08014__A1 _03252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06181__I _01612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12643__CLK net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06576__A1 _02078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10372__A2 _04962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09939_ _04579_ _04640_ _04641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09514__A1 u_cpu.rf_ram.memory\[33\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08317__A2 _03517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06328__A1 _01400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11901_ _00597_ net469 u_cpu.rf_ram.memory\[132\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11832_ _00528_ net478 u_cpu.rf_ram.memory\[138\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12023__CLK net495 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09817__A2 _04485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07828__A1 u_cpu.rf_ram.memory\[129\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11763_ _00459_ net491 u_cpu.rf_ram.memory\[141\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06187__S0 _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10714_ _05142_ _05176_ _05183_ _01139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11694_ _00398_ net329 u_cpu.rf_ram.memory\[56\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06500__B2 _02113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06351__I1 u_cpu.rf_ram.memory\[21\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12173__CLK net386 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08628__I0 _03566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10645_ _04820_ _05140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07056__A2 _02656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08253__A1 _03410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10576_ _02789_ _05098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10060__A1 _04411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12315_ _00995_ net528 u_cpu.cpu.ctrl.o_ibus_adr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xu_scanchain_local.scan_flop\[41\] u_scanchain_local.module_data_in\[40\] net553 u_arbiter.o_wb_cpu_adr\[3\]
+ net21 u_scanchain_local.module_data_in\[41\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_108_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08005__A1 _03266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12246_ _00929_ net272 u_cpu.rf_ram.memory\[32\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12177_ _00860_ net387 u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06567__A1 _01637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10363__A2 _04906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07915__I _03077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11128_ u_cpu.rf_ram.memory\[27\]\[0\] _05447_ _05448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09505__A1 _04244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08308__A2 _03514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11059_ u_cpu.rf_ram.memory\[87\]\[5\] _05396_ _05400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11312__A1 _04907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10115__A2 _04739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout365_I net366 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06975__B _01408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout532_I net534 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06266__I _01665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08270_ _03486_ _03487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_60_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08492__A1 _03604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07295__A2 _02833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07221_ _02740_ _02792_ _02794_ _00034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06893__I2 u_cpu.rf_ram.memory\[86\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09577__I _04311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07152_ _02712_ _02734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__11540__CLK net249 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08244__A1 _03421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12666__CLK net286 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06103_ _01595_ _01720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09992__A1 _04401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10051__B2 _04531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09992__B2 _04528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07083_ _01374_ _02675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_12_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06034_ _01650_ _01651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_82_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08547__A2 _03659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout104 net105 net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout115 net120 net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_47_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10354__A2 _04906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout126 net129 net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_138_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout137 net139 net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout148 net156 net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07985_ u_cpu.rf_ram.memory\[68\]\[6\] _03303_ _03308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout159 net161 net159 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_25_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09724_ _01438_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[13\] _04449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_47_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06936_ u_cpu.rf_ram_if.rtrig1 _02543_ _02544_ _02545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_28_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12046__CLK net495 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10106__A2 _04710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11303__A1 _02906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07358__I0 _02870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09655_ u_cpu.rf_ram.memory\[113\]\[1\] _04385_ _04387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06405__S1 _01908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06867_ _01760_ _02448_ _02457_ _02476_ _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_23_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08606_ _03666_ _03700_ _03702_ _00511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05818_ _01456_ _01460_ _01462_ u_arbiter.o_wb_cpu_adr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09586_ _04339_ _04340_ _00854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06798_ _01647_ _02399_ _02408_ _02409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06730__A1 _02322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08537_ _03588_ _03655_ _03657_ _00487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05749_ _01399_ _01400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12196__CLK net396 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06176__I _01632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08468_ _03600_ _03609_ _03616_ _00459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07286__A2 _02833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07419_ _02907_ _02925_ _02932_ _00094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_91_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08399_ _03571_ _00435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08391__I _02857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10430_ _04992_ _04997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07038__A2 _02603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10042__A1 _02605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09983__A1 _04468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08786__A2 _03801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10361_ _02545_ _02586_ _04953_ _04955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_30_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09983__B2 _04680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06636__I2 u_cpu.rf_ram.memory\[74\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06341__S0 _01583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12100_ _00783_ net437 u_cpu.rf_ram.memory\[121\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10593__A2 _05104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10292_ u_cpu.cpu.ctrl.o_ibus_adr\[3\] _04907_ _04910_ u_cpu.cpu.ctrl.o_ibus_adr\[4\]
+ _04914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_65_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09735__A1 _04452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08538__A2 _03656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12031_ _00714_ net312 u_cpu.rf_ram.memory\[91\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06549__A1 _01802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11257__I _05522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12539__CLK net293 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08566__I _03497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12864_ u_scanchain_local.data_out net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11815_ _00511_ net477 u_cpu.rf_ram.memory\[143\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11746_ _00003_ net252 u_cpu.rf_ram.rdata\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08474__A1 _03606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06086__I _01702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07277__A2 _02817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11563__CLK net341 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12689__CLK net234 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11677_ _00381_ net286 u_cpu.rf_ram.memory\[58\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10628_ u_arbiter.i_wb_cpu_rdt\[30\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[14\]
+ _05123_ _05128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07029__A2 _02633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10033__A1 _04402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10033__B2 _04509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08777__A2 _03802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout113_I net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10559_ u_cpu.rf_ram.memory\[96\]\[2\] _05088_ _05089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06627__I2 u_cpu.rf_ram.memory\[82\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06788__A1 _02392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06332__S0 _01826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06883__S1 _01707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09726__A1 _04439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08529__A2 _03647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12229_ _00912_ net361 u_cpu.cpu.immdec.imm30_25\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12069__CLK net282 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10336__A2 _04936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06689__C _01733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout482_I net483 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07201__A2 u_cpu.cpu.o_wdata0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07770_ _03060_ _03168_ _03170_ _00207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05763__A2 u_cpu.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06721_ _02039_ _02332_ _02333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08701__A2 _03748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09440_ u_cpu.rf_ram.memory\[122\]\[4\] _04230_ _04233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08476__I _03620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06652_ _02255_ _02264_ _02265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06712__A1 _01735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07380__I _02757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11906__CLK net471 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09371_ _02857_ _04190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11116__B _01394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06583_ _02189_ _02191_ _02193_ _02195_ _01784_ _02196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_80_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08322_ _03510_ _03514_ _03523_ _00406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout26_I net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07268__A2 _02818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08253_ _03410_ _03473_ _03476_ _00384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07204_ u_cpu.rf_ram.memory\[82\]\[7\] _02732_ _02779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08184_ _03419_ _03428_ _03435_ _00356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09965__A1 _02679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07135_ u_cpu.rf_ram_if.rcnt\[0\] _02717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08768__A2 _03287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07066_ u_cpu.rf_ram_if.rdata0\[2\] _02662_ _02664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07440__A2 _02942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06874__S1 _01693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06017_ _01633_ _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09193__A2 _04057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11436__CLK net327 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07968_ _03297_ _00278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05754__A2 _01388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09707_ u_arbiter.i_wb_cpu_rdt\[15\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\]
+ _01439_ _04432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06919_ _02527_ _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07899_ _03059_ _03252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09638_ _04374_ _04375_ _00871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11586__CLK net248 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09569_ u_arbiter.i_wb_cpu_rdt\[6\] _04326_ _04321_ u_arbiter.i_wb_cpu_dbus_dat\[6\]
+ _04327_ u_arbiter.i_wb_cpu_dbus_dat\[7\] _04328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_15_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11600_ _00304_ net244 u_cpu.rf_ram.memory\[65\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12580_ _01259_ net166 u_cpu.rf_ram.memory\[111\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11531_ _00235_ net489 u_cpu.rf_ram.memory\[139\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08208__A1 _03423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11462_ _00166_ net297 u_cpu.rf_ram.memory\[47\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06219__B1 _01829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09956__A1 u_cpu.cpu.immdec.imm24_20\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10413_ _04192_ u_cpu.rf_ram.memory\[2\]\[3\] _04983_ _04987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08759__A2 _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11393_ _00097_ net249 u_cpu.rf_ram.memory\[78\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10344_ _04944_ _01008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__12211__CLK net353 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07431__A2 _02940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09708__A1 _04431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06490__I0 u_cpu.rf_ram.memory\[40\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10275_ _04827_ _04895_ _04902_ _00981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12014_ _00697_ net411 u_cpu.rf_ram.memory\[36\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09184__A2 _04064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06617__S1 _01908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07195__A1 _02734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12361__CLK net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08931__A2 _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08497__S _03633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout490 net492 net490 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_24_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08296__I _03506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08695__A1 _03755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xserv_1_567 io_oeb[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_73_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09644__B1 _04329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08998__A2 _03946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout230_I net231 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11729_ _00433_ net128 u_cpu.rf_ram.memory\[9\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout328_I net336 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10006__A1 _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07422__A2 _02929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12704__CLK net239 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08940_ _02766_ _03912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07375__I _02751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09175__A2 _04058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08871_ u_cpu.rf_ram.memory\[130\]\[5\] _03863_ _03867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06608__S1 _01895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07186__A1 u_cpu.rf_ram.memory\[82\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07822_ _03179_ _03204_ _03206_ _00223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08922__A2 _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07753_ _03071_ _03154_ _03159_ _00201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06704_ _01904_ _02315_ _01679_ _02316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_38_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07489__A2 _02970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07684_ _03108_ _00183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09423_ u_cpu.rf_ram.memory\[112\]\[6\] _04217_ _04222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06635_ _01929_ _02247_ _01932_ _02248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09354_ _04150_ _04173_ _04179_ _00783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06566_ u_cpu.rf_ram.memory\[8\]\[4\] u_cpu.rf_ram.memory\[9\]\[4\] u_cpu.rf_ram.memory\[10\]\[4\]
+ u_cpu.rf_ram.memory\[11\]\[4\] _01574_ _01838_ _02179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_107_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08305_ _03512_ _03514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06449__B1 _02059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08989__A2 _03935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09285_ u_cpu.rf_ram.memory\[117\]\[3\] _04133_ _04135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06839__I2 u_cpu.rf_ram.memory\[22\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06497_ _01882_ _02110_ _02111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06544__S0 _01792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08236_ _03412_ _03461_ _03466_ _00377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12234__CLK net263 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08167_ _03423_ _03408_ _03424_ _00350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10548__A2 _05073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07118_ _02633_ _02703_ _02615_ _02605_ _02704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_109_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08098_ _03353_ _03370_ _03379_ _00326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07049_ _02650_ u_cpu.rf_ram_if.rdata1\[2\] _02653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10060_ _04411_ _04429_ _04490_ _04749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_66_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08913__A2 _03883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06924__A1 u_arbiter.i_wb_cpu_dbus_we vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10720__A2 _05177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06775__I1 u_cpu.rf_ram.memory\[33\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10962_ u_cpu.rf_ram.memory\[85\]\[1\] _05337_ _05339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08677__A1 _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12701_ u_cpu.rf_ram_if.wdata1_r\[5\] net233 u_cpu.rf_ram_if.wdata1_r\[4\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10484__A1 _02803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10893_ _05282_ _05290_ _05297_ _01204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08844__I _03846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12632_ _01311_ net59 u_cpu.rf_ram.memory\[25\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10087__I1 u_arbiter.i_wb_cpu_rdt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10087__S _01441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12563_ _01242_ net159 u_cpu.rf_ram.memory\[110\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10787__A2 _05219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11514_ _00218_ net320 u_cpu.rf_ram.memory\[119\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12494_ _01173_ net39 u_cpu.rf_ram.memory\[106\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09929__A1 _04397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11445_ _00149_ net325 u_cpu.rf_ram.memory\[43\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11601__CLK net243 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10539__A2 _05076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11376_ _00080_ net134 u_cpu.rf_ram.memory\[7\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10327_ _04934_ _01001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_84_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11751__CLK net479 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09157__A2 _04049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10258_ _04888_ _04891_ _04892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10011__I1 u_arbiter.i_wb_cpu_rdt\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08904__A2 _03886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09952__I1 u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10189_ u_arbiter.i_wb_cpu_dbus_adr\[5\] u_arbiter.i_wb_cpu_dbus_adr\[4\] _04849_
+ _04852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_78_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07963__I0 _02867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout180_I net183 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout278_I net279 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06539__I _01627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08668__A1 u_cpu.rf_ram.memory\[39\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout445_I net446 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06420_ _01772_ _02034_ _02035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09617__B1 _04359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12257__CLK net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07891__A2 _03245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06351_ u_cpu.rf_ram.memory\[20\]\[2\] u_cpu.rf_ram.memory\[21\]\[2\] u_cpu.rf_ram.memory\[22\]\[2\]
+ u_cpu.rf_ram.memory\[23\]\[2\] _01849_ _01965_ _01966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_37_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10778__A2 _05220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09070_ _03977_ _03991_ _03996_ _00681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06282_ u_cpu.rf_ram.memory\[96\]\[1\] u_cpu.rf_ram.memory\[97\]\[1\] u_cpu.rf_ram.memory\[98\]\[1\]
+ u_cpu.rf_ram.memory\[99\]\[1\] _01729_ _01641_ _01898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_124_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08021_ _03262_ _03324_ _03330_ _00298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09972_ _04465_ _04666_ _04672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_fanout93_I net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08923_ _02744_ _03899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07038__C _02578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08929__I _03895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08854_ _03830_ _03848_ _03856_ _00605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06906__A1 _02496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07805_ u_cpu.rf_ram.memory\[119\]\[4\] _03189_ _03194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08785_ _03761_ _03803_ _03811_ _00581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05997_ _01613_ _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_22_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06382__A2 _01995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07736_ u_cpu.rf_ram.memory\[16\]\[4\] _03146_ _03149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08659__A1 _03684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07667_ u_cpu.rf_ram.memory\[50\]\[6\] _03094_ _03099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09406_ _04211_ _00803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06618_ _01746_ _02230_ _02231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07882__A2 _03242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07598_ u_cpu.rf_ram.memory\[48\]\[1\] _03049_ _03051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06549_ _01802_ _02162_ _01805_ _02163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09337_ u_cpu.rf_ram.memory\[118\]\[5\] _04165_ _04169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06517__S0 _01741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10769__A2 _05162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09268_ _04068_ _04117_ _04124_ _00752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07634__A2 _03064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06437__A3 _02051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08219_ _02864_ u_cpu.rf_ram.memory\[5\]\[4\] _03451_ _03456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_5_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06117__C _01733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09199_ _02558_ _02594_ _04079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11230_ _02722_ _05243_ _05510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11774__CLK net512 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11161_ _05451_ _05465_ _05470_ _01299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_49_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10112_ _02684_ u_cpu.cpu.immdec.imm24_20\[0\] _04797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11092_ _05418_ _05421_ _05422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_49_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10043_ _02539_ _02624_ _04735_ _04736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__05972__B _01588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08839__I _03846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07570__A1 _03000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11994_ _00013_ net259 u_cpu.rf_ram_if.rdata0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10102__C _04511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10945_ _04190_ u_cpu.rf_ram.memory\[10\]\[2\] _05326_ _05329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07873__A2 _03233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10876_ u_cpu.rf_ram.memory\[108\]\[7\] _05269_ _05287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05884__A1 _01473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12615_ _01294_ net56 u_cpu.rf_ram.memory\[27\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06308__B _01782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06094__I _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12546_ _01225_ net116 u_cpu.rf_ram.memory\[10\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07625__A2 _03064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12477_ _01156_ net190 u_cpu.rf_ram.memory\[79\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07918__I _03080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11428_ _00132_ net333 u_cpu.rf_ram.memory\[51\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11185__A2 _05477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11359_ _00063_ net68 u_cpu.rf_ram.memory\[20\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05939__A2 _01557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout395_I net539 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05920_ _01524_ _01542_ _01543_ u_arbiter.o_wb_cpu_adr\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08749__I _03789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07653__I _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05851_ _01452_ _01489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10696__A1 _05144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout562_I net563 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07561__A1 u_cpu.rf_ram.memory\[41\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08570_ u_cpu.rf_ram.memory\[71\]\[4\] _03674_ _03679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05782_ u_arbiter.i_wb_cpu_ibus_adr\[0\] _01431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10448__A1 _04566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07521_ _02915_ _03000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_19_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09302__A2 _04143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07452_ _02953_ _02954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07864__A2 _03230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06911__I1 u_cpu.rf_ram.memory\[129\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06403_ u_cpu.rf_ram.memory\[120\]\[2\] u_cpu.rf_ram.memory\[121\]\[2\] u_cpu.rf_ram.memory\[122\]\[2\]
+ u_cpu.rf_ram.memory\[123\]\[2\] _01741_ _01905_ _02018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_50_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07383_ _02904_ _02893_ _02905_ _00085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_17_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09122_ _04026_ _03123_ _04027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06334_ u_cpu.rf_ram.memory\[132\]\[1\] u_cpu.rf_ram.memory\[133\]\[1\] u_cpu.rf_ram.memory\[134\]\[1\]
+ u_cpu.rf_ram.memory\[135\]\[1\] _01831_ _01832_ _01950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08813__A1 _03830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09053_ u_cpu.rf_ram.memory\[123\]\[5\] _03978_ _03985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10455__S _05004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06265_ _01691_ _01880_ _01695_ _01881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08004_ u_cpu.rf_ram.memory\[67\]\[5\] _03316_ _03320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06196_ _01812_ _01813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_89_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11176__A2 _05477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09955_ _04585_ _04655_ _04656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08906_ u_cpu.rf_ram.memory\[22\]\[3\] _03886_ _03888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09886_ _04249_ _04588_ _04595_ _00899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12422__CLK net363 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10687__A1 _05135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08837_ _03002_ _03814_ _03846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08768_ _03201_ _03287_ _03801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07719_ _01820_ _03136_ _03138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_2759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06107__A2 _01722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08699_ _03503_ _03759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12572__CLK net200 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08394__I _02860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10730_ _05137_ _05188_ _05193_ _01145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07855__A2 _03217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10661_ _05150_ _05151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09057__A1 _03986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06128__B _01744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05961__S1 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12400_ _01079_ net44 u_cpu.rf_ram.memory\[96\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08804__A1 _03824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10592_ _05053_ _05101_ _05108_ _01092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07607__A2 _03052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12331_ _01011_ net501 u_cpu.cpu.ctrl.o_ibus_adr\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12262_ _00945_ net491 u_arbiter.i_wb_cpu_dbus_adr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08407__I1 u_cpu.rf_ram.memory\[9\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11167__A2 _05466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11213_ _05500_ _05501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_135_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput6 net6 io_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_123_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12193_ _00876_ net403 u_cpu.rf_ram.memory\[113\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10914__A2 _05303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11144_ u_cpu.rf_ram.memory\[27\]\[5\] _05452_ _05459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09780__A2 _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06433__I3 u_cpu.rf_ram.memory\[79\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11075_ u_cpu.rf_ram.memory\[88\]\[3\] _05408_ _05410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08569__I _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[24\]_CLK net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07473__I _02966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10026_ _01440_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[7\] _04720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_114_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06346__A2 _01960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07543__A1 _02996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06310__C _01925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06089__I _01658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[39\]_CLK net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09296__A1 _03165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11977_ _00017_ net265 u_cpu.rf_ram_if.rdata1\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07846__A2 _03220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10928_ _05275_ _05314_ _05319_ _01217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05857__A1 _01489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout143_I net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09048__A1 _03980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10859_ _04816_ _05275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_125_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09843__I0 u_arbiter.i_wb_cpu_rdt\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout310_I net311 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12529_ _01208_ net276 u_cpu.rf_ram.memory\[84\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout408_I net412 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07648__I _03086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06050_ _01623_ _01667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.output_buffers\[3\] net34 u_scanchain_local.clk_out vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08023__A2 _03324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09220__A1 u_cpu.rf_ram.memory\[92\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10905__A2 _05302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12445__CLK net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09771__A2 _04493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout308 net311 net308 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_87_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout319 net320 net319 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_99_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06585__A2 _02197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07782__A1 u_cpu.rf_ram.memory\[40\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09740_ net8 _01433_ _04463_ _04464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06952_ _02559_ _02555_ _02557_ _02560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
.ends

