* NGSPICE file created from serv_1.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__sdffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__sdffq_1 D SE SI CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnq_1 D CLKN Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

.subckt serv_1 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_oeb[0] io_oeb[1] io_oeb[2]
+ io_oeb[3] io_oeb[4] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] vdd vss
XFILLER_41_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07909__I0 _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09523__A2 _04654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05903_ _02332_ u_cpu.cpu.mem_bytecnt\[1\] u_cpu.cpu.mem_bytecnt\[0\] _01409_ _02385_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09671_ _00125_ io_in[4] u_cpu.rf_ram.memory\[44\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06883_ u_cpu.rf_ram.memory\[60\]\[6\] _03002_ _03009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06337__A2 _02686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07534__A1 _03349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08622_ u_arbiter.i_wb_cpu_dbus_adr\[30\] _02445_ _04134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05834_ _02311_ u_cpu.cpu.immdec.imm31 _02317_ _02318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_55_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09287__A1 _04484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05765_ u_cpu.rf_ram.memory\[32\]\[7\] u_cpu.rf_ram.memory\[33\]\[7\] u_cpu.rf_ram.memory\[34\]\[7\]
+ u_cpu.rf_ram.memory\[35\]\[7\] _01623_ _01624_ _02250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08553_ _03547_ _04094_ _04098_ _00938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07504_ u_cpu.rf_ram.memory\[22\]\[6\] _03345_ _03358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08484_ _03782_ _04037_ _04046_ _03797_ _04047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_51_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07837__A2 _03541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05696_ _01541_ _02181_ _02182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[45\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05848__A1 _01369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07435_ _03161_ _03315_ _03317_ _00600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07366_ u_cpu.rf_ram.memory\[135\]\[3\] _03275_ _03279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09105_ u_cpu.rf_ram.memory\[106\]\[1\] _04419_ _04421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06317_ u_cpu.rf_ram.memory\[44\]\[2\] _02673_ _02676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07297_ _03167_ _03235_ _03240_ _00539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10417__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06273__A1 _02625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09036_ _04286_ _04379_ _04382_ _01137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06248_ u_cpu.rf_ram.memory\[78\]\[6\] _02628_ _02635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06179_ _02591_ _00070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08014__A2 _03648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05078__I _01398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05459__S0 _01680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10567__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06576__A2 _02834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09938_ _00392_ io_in[4] u_cpu.rf_ram.memory\[56\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09514__A2 _04654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09869_ _00323_ io_in[4] u_cpu.rf_ram.memory\[29\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06328__A2 _02673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07828__A2 _03541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10713_ _01142_ io_in[4] u_cpu.rf_ram.memory\[104\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06500__A2 _02791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10644_ _01073_ io_in[4] u_cpu.rf_ram.memory\[95\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10575_ _01005_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10097__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08253__A2 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09450__A1 _04482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06264__A1 _02497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08005__A2 u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[34\] u_arbiter.i_wb_cpu_rdt\[31\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[28\]
+ u_scanchain_local.clk u_scanchain_local.module_data_in\[34\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__07764__A1 _03359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06567__A2 _02823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11058_ _11058_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__09505__A2 _04644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06319__A2 _02673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07516__A1 _03349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10009_ _00455_ io_in[4] u_cpu.rf_ram.memory\[141\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[68\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05622__S0 _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09269__A1 _04484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05550_ _01399_ _02037_ _02038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08963__S _04331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05481_ u_cpu.rf_ram.memory\[28\]\[4\] u_cpu.rf_ram.memory\[29\]\[4\] u_cpu.rf_ram.memory\[30\]\[4\]
+ u_cpu.rf_ram.memory\[31\]\[4\] _01572_ _01574_ _01969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_20_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07220_ _03161_ _03196_ _03198_ _00504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08619__I1 u_arbiter.i_wb_cpu_dbus_adr\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07151_ _02599_ u_cpu.rf_ram.memory\[13\]\[7\] _03148_ _03156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09732__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08244__A2 _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06102_ _02482_ _02541_ _02542_ _00042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06255__A1 _02638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07082_ _02625_ _02832_ _03118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06033_ _02477_ _02487_ _02488_ _00027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07055__I0 _02587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09882__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08203__S _01436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06558__A2 _02823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07984_ _03553_ _03626_ _03633_ _00834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_47_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09723_ _00177_ io_in[4] u_cpu.rf_ram.memory\[50\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_101_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06935_ _02965_ _03031_ _03037_ _00380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08704__B1 _04175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09654_ _00108_ io_in[4] u_cpu.rf_ram.memory\[46\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06866_ _02967_ _02992_ _02999_ _00349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08180__A1 _03773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05613__S0 _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08605_ u_arbiter.i_wb_cpu_dbus_adr\[23\] u_arbiter.i_wb_cpu_dbus_adr\[22\] _04115_
+ _04125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05817_ _02295_ _02297_ _02299_ _02301_ _01404_ _02302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_09585_ _00039_ io_in[4] u_cpu.rf_ram.memory\[21\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06797_ _02491_ _02959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08307__I0 u_arbiter.i_wb_cpu_rdt\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06730__A2 _02914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08536_ u_cpu.rf_ram.memory\[32\]\[4\] _04084_ _04089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05748_ _01542_ _02232_ _01417_ _02233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_23_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05679_ _02158_ _02160_ _02162_ _02164_ _01628_ _02165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_08467_ _03890_ _03790_ _04031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05297__A2 _01786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06494__A1 _02769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07418_ u_cpu.rf_ram.memory\[132\]\[2\] _03305_ _03308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08398_ _03743_ _03786_ _03828_ _03831_ _03904_ _03970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_104_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07349_ _03165_ _03265_ _03269_ _00562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09432__A1 _04482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10360_ _00793_ io_in[4] u_cpu.rf_ram.memory\[8\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07994__A1 _03545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09019_ u_cpu.rf_ram.memory\[103\]\[3\] _04369_ _04373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10291_ _00724_ io_in[4] u_cpu.rf_ram.memory\[90\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06549__A2 _02812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07746__A1 _01428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09499__A1 _04478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09605__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08171__A1 _03754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05524__A3 _02011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06721__A2 _02914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09755__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06485__A1 u_arbiter.i_wb_cpu_ack vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05288__A2 _01778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10732__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10627_ _01056_ io_in[4] u_cpu.rf_ram.memory\[97\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08226__A2 _03798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[2\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06237__A1 _02482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05220__B _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10558_ _00988_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06788__A2 _02944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10489_ _00922_ io_in[4] u_cpu.cpu.immdec.imm19_12_20\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10882__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07737__A1 _01408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08250__C _03835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10112__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04981_ _01443_ _01486_ _01488_ _01489_ u_arbiter.o_wb_cpu_adr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_110_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06960__A2 _03051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06720_ _02738_ _02914_ _02915_ _00287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06651_ u_cpu.rf_ram.memory\[76\]\[2\] _02874_ _02877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06712__A2 _02904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05602_ _02082_ _02084_ _02086_ _02088_ _01628_ _02089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_18_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10262__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05071__S1 _01557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09370_ _04569_ _04573_ _04574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06582_ _02746_ _02834_ _02838_ _00226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05920__B1 _01381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05533_ _02014_ _02016_ _02018_ _02020_ _01426_ _02021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_08321_ _03742_ _03900_ _03901_ _03902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_75_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08465__A2 _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06476__A1 _01372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08252_ _03740_ _03844_ _03845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05279__A2 _01760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05464_ _01684_ _01952_ _01418_ _01953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07203_ u_cpu.rf_ram.memory\[71\]\[2\] _03186_ _03189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08183_ _03763_ _03782_ _03783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09414__A1 _04482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05395_ u_cpu.rf_ram.memory\[24\]\[3\] u_cpu.rf_ram.memory\[25\]\[3\] u_cpu.rf_ram.memory\[26\]\[3\]
+ u_cpu.rf_ram.memory\[27\]\[3\] _01578_ _01580_ _01884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_118_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07134_ u_cpu.rf_ram.memory\[140\]\[7\] _03139_ _03147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07976__A1 _03545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06779__A2 _02944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07065_ _02577_ _02727_ _03109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07836__I _02506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06016_ u_cpu.cpu.immdec.imm11_7\[4\] _02457_ _02472_ _02473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_82_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05451__A2 _01939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08776__I0 _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09628__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05203__A2 _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07967_ u_cpu.rf_ram.memory\[115\]\[7\] _03616_ _03624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06951__A2 _03041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09706_ _00160_ io_in[4] u_cpu.rf_ram.memory\[48\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06918_ _02596_ u_cpu.rf_ram.memory\[5\]\[6\] _03021_ _03028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10605__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08153__A1 _01436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07898_ _02577_ _02706_ _03586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09637_ _00091_ io_in[4] u_cpu.rf_ram.memory\[78\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06849_ u_cpu.rf_ram.memory\[62\]\[7\] _02982_ _02990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09778__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06703__A2 _02904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09568_ _04687_ _01364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10755__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08519_ u_arbiter.i_wb_cpu_rdt\[31\] u_arbiter.i_wb_cpu_rdt\[15\] _01437_ _04078_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_90_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09499_ _04478_ _04644_ _04649_ _01333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08456__A2 _04016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06219__A1 _02492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10412_ _00845_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10343_ _00776_ io_in[4] u_cpu.rf_ram.memory\[118\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10274_ _00707_ io_in[4] u_cpu.cpu.state.o_cnt_r\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10135__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07719__A1 _03351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08778__S _04217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07195__A2 _03176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08392__A1 _03812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08519__I0 u_arbiter.i_wb_cpu_rdt\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06942__A2 _03041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10285__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05130__A1 _01589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07258__I0 _02587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05681__A2 _02138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05180_ _01553_ _01671_ _01565_ _01672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_122_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07958__A1 _03545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08080__B1 _03654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06630__A1 _02738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08870_ _04288_ _04282_ _04289_ _01064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10628__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05176__I _01548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07186__A2 _03176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07821_ _03540_ _03541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06933__A2 _03031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09920__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07752_ _03347_ _03500_ _03502_ _00733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_04964_ u_arbiter.i_wb_cpu_dbus_adr\[11\] _01457_ _01477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__04944__A1 _01445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05292__S1 _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08135__A1 _03551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06703_ u_cpu.rf_ram.memory\[68\]\[1\] _02904_ _02906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10778__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07683_ u_cpu.cpu.state.o_cnt_r\[3\] _03458_ _03459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04895_ _01419_ _01420_ _01421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08686__A2 _04155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09422_ _04472_ _04605_ _04607_ _01298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_92_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06634_ _02744_ _02864_ _02867_ _00249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09353_ _04478_ _04556_ _04561_ _01275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06565_ _02748_ _02823_ _02828_ _00219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10008__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08304_ _03553_ _03879_ _03886_ _00901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05516_ _01398_ _02003_ _02004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09284_ u_cpu.rf_ram.memory\[110\]\[6\] _04516_ _04523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06496_ _01681_ _02786_ _02789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_138_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07110__A2 _03129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05121__A1 _01609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08235_ u_arbiter.i_wb_cpu_rdt\[12\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[12\]
+ _01435_ _03830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05447_ _01667_ _01935_ _01936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05672__A2 _02157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08166_ _01435_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[14\] _03766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05378_ _01858_ _01867_ _01868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10158__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07117_ _02969_ _03129_ _03137_ _00462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08097_ u_arbiter.i_wb_cpu_rdt\[23\] _03653_ _03654_ u_arbiter.i_wb_cpu_dbus_dat\[23\]
+ _03714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_106_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07048_ _02577_ _02695_ _03100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08749__I0 _02573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05086__I _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07177__A2 _03159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08374__A1 _03797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08999_ u_cpu.rf_ram.memory\[102\]\[2\] _04359_ _04362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06924__A2 _03031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05283__S1 _01681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04935__A1 _01445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10961_ _10961_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_43_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10892_ _01321_ io_in[4] u_cpu.rf_ram.memory\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06860__A1 _02961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05663__A2 _02148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06612__A1 _02738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10326_ _00759_ io_in[4] u_cpu.rf_ram.memory\[117\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09943__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10257_ _00690_ io_in[4] u_cpu.rf_ram.memory\[37\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07168__A2 _03159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08365__A1 _03773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10188_ _00634_ io_in[4] u_cpu.rf_ram.memory\[128\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10920__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05274__S1 _01668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08668__A2 _04155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07340__A2 _02832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07479__I0 _02596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06350_ _02521_ _02637_ _02695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_72_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08971__S _04331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09093__A2 _04409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05301_ u_cpu.rf_ram.memory\[20\]\[2\] u_cpu.rf_ram.memory\[21\]\[2\] u_cpu.rf_ram.memory\[22\]\[2\]
+ u_cpu.rf_ram.memory\[23\]\[2\] _01572_ _01574_ _01791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10300__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06281_ u_cpu.rf_ram.memory\[46\]\[3\] _02651_ _02655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05232_ _01609_ _01722_ _01723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08020_ u_arbiter.i_wb_cpu_dbus_dat\[1\] _03650_ _03659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06851__A1 _02660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05163_ _01614_ _01653_ _01654_ _01655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_7_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10952__D u_cpu.rf_ram_if.wdata1_r\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10450__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09971_ _00425_ io_in[4] u_cpu.rf_ram.memory\[52\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05094_ u_cpu.rf_ram.memory\[24\]\[0\] u_cpu.rf_ram.memory\[25\]\[0\] u_cpu.rf_ram.memory\[26\]\[0\]
+ u_cpu.rf_ram.memory\[27\]\[0\] _01578_ _01580_ _01586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08922_ _01437_ _04319_ _04320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07159__A2 _03159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08853_ u_cpu.rf_ram.memory\[97\]\[6\] _04271_ _04278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07804_ _03343_ _03530_ _03531_ _00756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05265__S1 _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04917__A1 _01437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08784_ u_cpu.rf_ram.memory\[93\]\[0\] _04227_ _04228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05996_ u_cpu.cpu.bufreg.lsb\[1\] _02455_ _02332_ u_arbiter.i_wb_cpu_dbus_sel\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_73_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07735_ _02328_ _03489_ _03490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_38_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05590__A1 _01645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04947_ _01461_ _01462_ _01463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07666_ _03355_ _03442_ _03448_ _00700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_04878_ _01377_ _01387_ _01403_ _01404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07331__A2 _03255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09405_ u_cpu.rf_ram.memory\[27\]\[2\] _04595_ _04598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06617_ u_cpu.rf_ram.memory\[77\]\[3\] _02854_ _02858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05342__A1 _01645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07597_ u_cpu.rf_ram.memory\[124\]\[7\] _03402_ _03410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09336_ u_cpu.rf_ram.memory\[87\]\[5\] _04546_ _04552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06548_ _02750_ _02812_ _02818_ _00212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09816__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07095__A1 _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09267_ _04482_ _04506_ _04513_ _01237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06479_ u_arbiter.i_wb_cpu_dbus_dat\[0\] u_arbiter.i_wb_cpu_dbus_dat\[1\] u_arbiter.i_wb_cpu_dbus_dat\[2\]
+ u_arbiter.i_wb_cpu_dbus_dat\[3\] _02775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_138_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08218_ _03815_ _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05645__A2 _02130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06842__A1 _02961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07890__I0 _02590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09198_ _04472_ _04470_ _04473_ _01208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08149_ _03748_ _03749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09966__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07398__A2 _03295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10943__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10111_ _00557_ io_in[4] u_cpu.rf_ram.memory\[49\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11091_ _11091_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08347__A1 _03831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10042_ _00488_ io_in[4] u_cpu.rf_ram.memory\[73\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08898__A2 _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04869__B _01387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04908__A1 u_arbiter.i_wb_cpu_ibus_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07570__A2 _03392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05581__A1 _01601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10944_ _01364_ io_in[4] u_cpu.rf_ram_if.rgnt vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07322__A2 _02684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10323__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05333__A1 _01594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10875_ _01304_ io_in[4] u_cpu.rf_ram.memory\[26\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09075__A2 _04399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05212__C _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[64\] u_scanchain_local.module_data_in\[63\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[26\] u_scanchain_local.clk u_scanchain_local.module_data_in\[64\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__08804__B _03788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10473__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06833__A1 _02625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05636__A2 _02122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07389__A2 _03285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10309_ _00742_ io_in[4] u_cpu.rf_ram.memory\[35\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05495__S1 _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08338__A1 u_cpu.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08889__A2 _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05850_ u_cpu.cpu.bne_or_bge _02333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_120_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07561__A2 _03382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05781_ u_cpu.rf_ram.memory\[120\]\[7\] u_cpu.rf_ram.memory\[121\]\[7\] u_cpu.rf_ram.memory\[122\]\[7\]
+ u_cpu.rf_ram.memory\[123\]\[7\] _01646_ _01603_ _02266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_35_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05572__A1 _01542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07520_ _03353_ _03362_ _03367_ _00635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09839__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08510__A1 _01437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07313__A2 _03245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05324__A1 _01589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07451_ _03157_ _03325_ _03326_ _00607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06402_ u_cpu.rf_ram.memory\[48\]\[6\] _02718_ _02725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10816__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07382_ u_cpu.rf_ram.memory\[134\]\[2\] _03285_ _03288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09121_ u_cpu.rf_ram.memory\[107\]\[0\] _04429_ _04430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06333_ _02685_ _02686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09989__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09052_ _04284_ _04389_ _04391_ _01144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06264_ _02497_ _02641_ _02645_ _00101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05627__A2 _02113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06824__A1 _02961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05183__S0 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08003_ u_cpu.rf_ram.memory\[33\]\[7\] _03636_ _03644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08433__C _03755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05215_ u_cpu.rf_ram.memory\[16\]\[1\] u_cpu.rf_ram.memory\[17\]\[1\] u_cpu.rf_ram.memory\[18\]\[1\]
+ u_cpu.rf_ram.memory\[19\]\[1\] _01578_ _01580_ _01706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_06195_ _02573_ u_cpu.rf_ram.memory\[7\]\[0\] _02603_ _02604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05146_ _01636_ _01637_ _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05077_ _01552_ _01559_ _01561_ _01566_ _01568_ _01569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_09954_ _00408_ io_in[4] u_cpu.rf_ram.memory\[54\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05486__S1 _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08329__A1 _03767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08905_ u_cpu.rf_ram.memory\[96\]\[1\] _04309_ _04311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09885_ _00339_ io_in[4] u_cpu.rf_ram.memory\[62\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07001__A1 _02959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08836_ _03740_ _03741_ _04267_ _04268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07552__A2 _03382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10346__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05563__A1 _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08767_ _04218_ _01032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_122_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05979_ _01372_ _02394_ _02441_ _02443_ _02444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_73_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07718_ u_cpu.rf_ram.memory\[90\]\[3\] _03475_ _03479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08698_ u_cpu.cpu.ctrl.o_ibus_adr\[19\] _04173_ _04175_ u_cpu.cpu.ctrl.o_ibus_adr\[20\]
+ _04179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_53_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08501__A1 _03742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07304__A2 _02832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07649_ u_cpu.rf_ram.memory\[37\]\[6\] _03432_ _03439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05315__A1 _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10496__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05866__A2 _02348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05313__B _01564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10660_ _01089_ io_in[4] u_cpu.rf_ram.memory\[28\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09057__A2 _04389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09319_ _04480_ _04536_ _04542_ _01260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10591_ _01021_ io_in[4] u_cpu.rf_ram.memory\[109\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08804__A2 _03818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08624__B _02445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05618__A2 _02104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06815__A1 _02684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05477__S1 _01574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07240__A1 _03163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07791__A2 _03520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11074_ _11074_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_62_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10025_ _00471_ io_in[4] u_cpu.rf_ram.memory\[13\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07543__A2 _03372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05554__A1 _02032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10839__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09296__A2 _04526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05306__A1 _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10927_ _01355_ io_in[4] u_cpu.rf_ram.memory\[23\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05857__A2 u_cpu.cpu.state.o_cnt_r\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10858_ _01287_ io_in[4] u_cpu.cpu.ctrl.i_iscomp vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10789_ _01218_ io_in[4] u_cpu.rf_ram.memory\[59\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06282__A2 _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10219__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08559__A1 _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05000_ u_cpu.cpu.ctrl.o_ibus_adr\[20\] _01498_ _01503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09220__A2 _04487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05893__B _01373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05468__S1 _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07782__A2 _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10369__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06951_ _02963_ _03041_ _03046_ _00387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05902_ u_cpu.cpu.mem_if.signbit _02384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_39_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09670_ _00124_ io_in[4] u_cpu.rf_ram.memory\[44\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06882_ _02965_ _03002_ _03008_ _00356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09661__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07534__A2 _03372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08621_ u_arbiter.i_wb_cpu_dbus_adr\[31\] _04133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_94_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05833_ _01369_ _01372_ _01374_ _02317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08552_ u_cpu.rf_ram.memory\[31\]\[3\] _04094_ _04098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05764_ _01597_ _02248_ _02249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09287__A2 _04516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07503_ _02511_ _03357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_78_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08483_ _04038_ _04039_ _03782_ _04045_ _04046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_05695_ u_cpu.rf_ram.memory\[112\]\[6\] u_cpu.rf_ram.memory\[113\]\[6\] u_cpu.rf_ram.memory\[114\]\[6\]
+ u_cpu.rf_ram.memory\[115\]\[6\] _01619_ _01620_ _02181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__05848__A2 _02309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07434_ u_cpu.rf_ram.memory\[131\]\[1\] _03315_ _03317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09039__A2 _04379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07365_ _03163_ _03275_ _03278_ _00569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09104_ _04280_ _04419_ _04420_ _01167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07839__I _02511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06316_ _02487_ _02673_ _02675_ _00123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05787__C _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07296_ u_cpu.rf_ram.memory\[39\]\[4\] _03235_ _03240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09035_ u_cpu.rf_ram.memory\[104\]\[2\] _04379_ _04382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06273__A2 _02639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06247_ _02507_ _02628_ _02634_ _00095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06178_ _02590_ u_cpu.rf_ram.memory\[1\]\[4\] _02578_ _02591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_104_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07222__A1 _03163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05129_ u_cpu.rf_ram.memory\[36\]\[0\] u_cpu.rf_ram.memory\[37\]\[0\] u_cpu.rf_ram.memory\[38\]\[0\]
+ u_cpu.rf_ram.memory\[39\]\[0\] _01619_ _01620_ _01621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__05459__S1 _01681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07773__A2 _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09937_ _00391_ io_in[4] u_cpu.rf_ram.memory\[56\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05784__A1 _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05308__B _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09868_ _00322_ io_in[4] u_cpu.rf_ram.memory\[29\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08722__A1 _02343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07525__A2 _03362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08819_ _03812_ _04252_ _04253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_45_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09799_ _00253_ io_in[4] u_cpu.rf_ram.memory\[74\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09278__A2 _04516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07289__A1 _03157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10712_ _01141_ io_in[4] u_cpu.rf_ram.memory\[104\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05839__A2 _02320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05395__S0 _01578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10643_ _01072_ io_in[4] u_cpu.rf_ram.memory\[95\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08789__A1 _03545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05147__S0 _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10574_ _01004_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09450__A2 _04615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06264__A2 _02641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07461__A1 _03169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10511__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[27\] u_arbiter.i_wb_cpu_rdt\[24\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[21\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_123_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09684__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07764__A2 _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05775__A1 _01636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11057_ _11057_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_114_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10661__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07516__A2 _03362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10008_ _00454_ io_in[4] u_cpu.rf_ram.memory\[142\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05622__S1 _01668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09269__A2 _04506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05480_ _01562_ _01967_ _01582_ _01968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_60_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05386__S0 _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08229__B1 _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08264__B _03855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10041__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07150_ _03155_ _00477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09441__A2 _04615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06101_ u_cpu.rf_ram.memory\[81\]\[0\] _02541_ _02542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06255__A2 _02639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07081_ _03117_ _00446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06032_ u_cpu.rf_ram.memory\[82\]\[1\] _02477_ _02488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10191__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07204__A1 _03163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07755__A2 _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05766__A1 _01645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07983_ u_cpu.rf_ram.memory\[116\]\[6\] _03626_ _03633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05310__S0 _01590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09722_ _00176_ io_in[4] u_cpu.rf_ram.memory\[50\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_101_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06934_ u_cpu.rf_ram.memory\[58\]\[5\] _03031_ _03037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[12\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07507__A2 _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09653_ _00107_ io_in[4] u_cpu.rf_ram.memory\[46\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05518__A1 _01645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06865_ u_cpu.rf_ram.memory\[61\]\[6\] _02992_ _02999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08180__A2 _03755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08604_ _04124_ _00963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05816_ _01684_ _02300_ _01418_ _02301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05613__S1 _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09584_ _00038_ io_in[4] u_cpu.rf_ram.memory\[21\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06796_ _02957_ _02955_ _02958_ _00320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08307__I1 u_arbiter.i_wb_cpu_rdt\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08535_ _03547_ _04084_ _04088_ _00930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05747_ u_cpu.rf_ram.memory\[24\]\[7\] u_cpu.rf_ram.memory\[25\]\[7\] u_cpu.rf_ram.memory\[26\]\[7\]
+ u_cpu.rf_ram.memory\[27\]\[7\] _01578_ _01580_ _02232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_24_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08466_ _03835_ _03988_ _04030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05678_ _01645_ _02163_ _01626_ _02164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07417_ _03161_ _03305_ _03307_ _00592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06494__A2 _02783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08397_ _03762_ _03891_ _03894_ _03969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[23\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07348_ u_cpu.rf_ram.memory\[136\]\[3\] _03265_ _03269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05129__S0 _01619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09432__A2 _04605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10534__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06246__A2 _02628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07443__A1 _03169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07279_ _03167_ _03225_ _03230_ _00531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07994__A2 _03636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09018_ _04286_ _04369_ _04372_ _01129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10290_ _00723_ io_in[4] u_cpu.rf_ram.memory\[90\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[38\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10684__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05757__A1 _01601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05301__S0 _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09499__A2 _04644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05509__A1 _01594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04980__A2 _01442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08171__A2 _03755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10064__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06485__A2 _01442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07682__A1 _01428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10626_ _01055_ io_in[4] u_cpu.rf_ram.memory\[97\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09423__A2 _04605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06237__A2 _02628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10557_ _00987_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07985__A2 _03626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05540__S0 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05996__A1 u_cpu.cpu.bufreg.lsb\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10488_ _00921_ io_in[4] u_cpu.cpu.immdec.imm19_12_20\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07737__A2 _02332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[35\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05748__A1 _01542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11109_ io_oeb[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_96_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04980_ u_arbiter.i_wb_cpu_dbus_adr\[15\] _01442_ _01489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08698__B1 _04175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04971__A2 _01442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10407__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06650_ _02742_ _02874_ _02876_ _00256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05601_ _01594_ _02087_ _01626_ _02088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06581_ u_cpu.rf_ram.memory\[129\]\[3\] _02834_ _02838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05920__A1 _01374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08320_ _03741_ _03831_ _03901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05532_ _01614_ _02019_ _01654_ _02020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_33_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10557__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06476__A2 _02332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08251_ _03767_ _03774_ _03801_ _03843_ _03844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_32_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05279__A3 _01769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05463_ u_cpu.rf_ram.memory\[132\]\[3\] u_cpu.rf_ram.memory\[133\]\[3\] u_cpu.rf_ram.memory\[134\]\[3\]
+ u_cpu.rf_ram.memory\[135\]\[3\] _01687_ _01688_ _01952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_123_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07202_ _03161_ _03186_ _03188_ _00496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08182_ _03774_ _03781_ _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05394_ _01570_ _01882_ _01883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09414__A2 _04595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06228__A2 _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07133_ _02967_ _03139_ _03146_ _00469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07425__A1 _03169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07976__A2 _03626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07064_ _03108_ _00438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05987__A1 u_arbiter.i_wb_cpu_ibus_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05531__S0 _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09178__A1 _04284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06015_ _02471_ _02472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_47_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05739__A1 _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06400__A2 _02718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07966_ _03553_ _03616_ _03623_ _00826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09705_ _00159_ io_in[4] u_cpu.rf_ram.memory\[48\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06917_ _03027_ _00372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_74_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08689__B1 _04157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07897_ _03585_ _00795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10087__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09636_ _00090_ io_in[4] u_cpu.rf_ram.memory\[78\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06468__I _01435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06848_ _02967_ _02982_ _02989_ _00341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05598__S0 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09567_ _01429_ u_cpu.rf_ram_if.rreq_r _04687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_130_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05911__A1 u_cpu.cpu.immdec.imm31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06779_ u_cpu.rf_ram.memory\[64\]\[3\] _02944_ _02948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08518_ _03835_ _03988_ _03902_ _03899_ _04077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_12_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09498_ u_cpu.rf_ram.memory\[98\]\[4\] _04644_ _04649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07664__A1 _03353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08449_ u_cpu.cpu.immdec.imm19_12_20\[1\] _03798_ _04016_ _04017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05770__S0 _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09405__A2 _04595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06219__A2 _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10411_ _00844_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07967__A2 _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[58\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10342_ _00775_ io_in[4] u_cpu.rf_ram.memory\[118\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08351__C _03826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10273_ _00706_ io_in[4] u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07719__A2 _03475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08916__A1 _04294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08519__I1 u_arbiter.i_wb_cpu_rdt\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__04953__A2 _01457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09722__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09341__A1 _04484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05589__S0 _01623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09872__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05761__S0 _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10609_ _01038_ io_in[4] u_cpu.rf_ram.memory\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07407__A1 _03169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05681__A3 _02147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07958__A2 _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08080__A1 u_arbiter.i_wb_cpu_rdt\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06630__A2 _02864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08969__S _04331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07820_ _02810_ _02821_ _03540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09373__B u_cpu.cpu.genblk3.csr.o_new_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07751_ u_cpu.rf_ram.memory\[92\]\[1\] _03500_ _03502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04963_ _01470_ _01461_ _01462_ _01475_ _01476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_65_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08135__A2 _03731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06702_ _02738_ _02904_ _02905_ _00279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_93_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07682_ _01428_ _02311_ _03458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06146__A1 _02497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04894_ u_cpu.cpu.immdec.imm24_20\[3\] _01388_ _01420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05192__I _01667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09421_ u_cpu.rf_ram.memory\[26\]\[1\] _04605_ _04607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06633_ u_cpu.rf_ram.memory\[74\]\[2\] _02864_ _02867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09352_ u_cpu.rf_ram.memory\[88\]\[4\] _04556_ _04561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06564_ u_cpu.rf_ram.memory\[119\]\[4\] _02823_ _02828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08303_ u_cpu.rf_ram.memory\[114\]\[6\] _03879_ _03886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05515_ u_cpu.rf_ram.memory\[124\]\[4\] u_cpu.rf_ram.memory\[125\]\[4\] u_cpu.rf_ram.memory\[126\]\[4\]
+ u_cpu.rf_ram.memory\[127\]\[4\] _01545_ _01642_ _02003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07646__A1 _03353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06449__A2 _02740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09283_ _04480_ _04516_ _04522_ _01244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06495_ _02788_ _00189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08234_ _03763_ _03790_ _03818_ _03827_ _03828_ _03802_ _03829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_05446_ u_cpu.rf_ram.memory\[64\]\[3\] u_cpu.rf_ram.memory\[65\]\[3\] u_cpu.rf_ram.memory\[66\]\[3\]
+ u_cpu.rf_ram.memory\[67\]\[3\] _01571_ _01668_ _01935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__05121__A2 _01612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05752__S0 _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09399__A1 _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08165_ _03757_ _03759_ _03764_ _03765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_101_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05377_ _01860_ _01862_ _01864_ _01866_ _01404_ _01867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__08452__B _04016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07949__A2 _03606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07116_ u_cpu.rf_ram.memory\[141\]\[7\] _03129_ _03137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08096_ u_arbiter.i_wb_cpu_dbus_dat\[24\] _03683_ _03713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06621__A2 _02854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07047_ _02969_ _03091_ _03099_ _00430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09745__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09571__A1 _02783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06385__A1 _02512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08998_ _04284_ _04359_ _04361_ _01120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07949_ u_cpu.rf_ram.memory\[122\]\[7\] _03606_ _03614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10722__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08126__A2 _03731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09323__A1 _04484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[1\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10960_ _10960_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_29_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06137__A1 _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09895__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09619_ _00073_ io_in[4] u_cpu.rf_ram.memory\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10891_ _01320_ io_in[4] u_cpu.rf_ram.memory\[24\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10872__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05743__S0 _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10102__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06860__A2 _02992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10325_ _00758_ io_in[4] u_cpu.rf_ram.memory\[117\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06612__A2 _02854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10252__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05966__A4 u_cpu.cpu.state.o_cnt_r\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10256_ _00689_ io_in[4] u_cpu.rf_ram.memory\[37\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08365__A2 _03767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09562__A1 _04155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10187_ _00633_ io_in[4] u_cpu.rf_ram.memory\[128\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04926__A2 _01443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06128__A1 _02502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07876__A1 _03551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06679__A2 _02884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07628__A1 _03353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05300_ _01783_ _01785_ _01787_ _01789_ _01568_ _01790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__09618__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06280_ _02492_ _02651_ _02654_ _00108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05734__S0 _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05231_ u_cpu.rf_ram.memory\[40\]\[1\] u_cpu.rf_ram.memory\[41\]\[1\] u_cpu.rf_ram.memory\[42\]\[1\]
+ u_cpu.rf_ram.memory\[43\]\[1\] _01610_ _01611_ _01722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_128_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06851__A2 _02684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04862__A1 u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05162_ _01564_ _01654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09768__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07800__A1 _03359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09970_ _00424_ io_in[4] u_cpu.rf_ram.memory\[52\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06603__A2 _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05093_ _01570_ _01584_ _01585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05257__I3 u_cpu.rf_ram.memory\[119\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08921_ u_arbiter.i_wb_cpu_ack u_arbiter.o_wb_cpu_adr\[1\] _04319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10745__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09553__A1 _04478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08356__A2 _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08852_ _03551_ _04271_ _04277_ _01058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07803_ u_cpu.rf_ram.memory\[117\]\[0\] _03530_ _03531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08783_ _04226_ _04227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05995_ u_cpu.cpu.bufreg.lsb\[0\] u_cpu.cpu.bne_or_bge _02455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08108__A2 _03676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09305__A1 _04484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07734_ _02325_ _03487_ _03489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_04946_ u_cpu.cpu.ctrl.o_ibus_adr\[7\] u_cpu.cpu.ctrl.o_ibus_adr\[6\] u_cpu.cpu.ctrl.o_ibus_adr\[5\]
+ _01451_ _01462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__10895__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05590__A2 _02076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07665_ u_cpu.rf_ram.memory\[36\]\[5\] _03442_ _03448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06914__I0 _02590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04877_ _01368_ _01403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08447__B _02767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09404_ _04472_ _04595_ _04597_ _01290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06616_ _02744_ _02854_ _02857_ _00241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07596_ _03357_ _03402_ _03409_ _00669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10125__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09335_ _04478_ _04546_ _04551_ _01267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06547_ u_cpu.rf_ram.memory\[40\]\[5\] _02812_ _02818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08292__A1 _03539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09266_ u_cpu.rf_ram.memory\[85\]\[6\] _04506_ _04513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07095__A2 _03119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06478_ _02772_ _02773_ _02774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05725__S0 _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08217_ _03796_ _03811_ _03815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05429_ u_cpu.rf_ram.memory\[120\]\[3\] u_cpu.rf_ram.memory\[121\]\[3\] u_cpu.rf_ram.memory\[122\]\[3\]
+ u_cpu.rf_ram.memory\[123\]\[3\] _01646_ _01603_ _01918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09197_ u_cpu.rf_ram.memory\[84\]\[1\] _04470_ _04473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06842__A2 _02982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10275__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08148_ _03745_ _03747_ _03748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_14_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08079_ _03701_ _03702_ _00860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05097__I _01397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10110_ _00556_ io_in[4] u_cpu.rf_ram.memory\[49\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11090_ _11090_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_96_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08347__A2 _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10041_ _00487_ io_in[4] u_cpu.rf_ram.memory\[73\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06358__A1 _02492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05825__I u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04869__C _01368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04908__A2 _01431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05581__A2 _02067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07858__A1 _03551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10943_ _01363_ io_in[4] u_cpu.rf_ram_if.rdata0\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10874_ _01303_ io_in[4] u_cpu.rf_ram.memory\[26\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10618__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08871__I _02501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08283__A1 _03762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07086__A2 _03119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05716__S0 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_scanchain_local.scan_flop\[57\] u_scanchain_local.module_data_in\[56\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[19\] u_scanchain_local.clk u_scanchain_local.module_data_in\[57\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__06833__A2 _02684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09910__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04904__I io_in[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10768__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10308_ _00741_ io_in[4] u_cpu.rf_ram.memory\[35\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09535__A1 _04478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08338__A2 _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10239_ _00008_ io_in[4] u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06349__A1 _02517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07010__A2 _03071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05021__A1 _01445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05780_ _01589_ _02264_ _02265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05411__I3 u_cpu.rf_ram.memory\[39\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07149__I0 _02596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05572__A2 _02058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10148__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07450_ u_cpu.rf_ram.memory\[130\]\[0\] _03325_ _03326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05324__A2 _01813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06521__A1 _02742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06401_ _02507_ _02718_ _02724_ _00159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07381_ _03161_ _03285_ _03287_ _00576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05875__A3 _02356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10298__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09120_ _04428_ _04429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06332_ _02682_ _02684_ _02685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08274__A1 _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05707__S0 _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09051_ u_cpu.rf_ram.memory\[99\]\[1\] _04389_ _04391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09590__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06263_ u_cpu.rf_ram.memory\[42\]\[3\] _02641_ _02645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06824__A2 _02972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05183__S1 _01549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08002_ _03553_ _03636_ _03643_ _00842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05214_ _01570_ _01704_ _01705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08026__A1 _03648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06194_ _02577_ _02602_ _02603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05145_ u_cpu.rf_ram.memory\[100\]\[0\] u_cpu.rf_ram.memory\[101\]\[0\] u_cpu.rf_ram.memory\[102\]\[0\]
+ u_cpu.rf_ram.memory\[103\]\[0\] _01598_ _01573_ _01637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_116_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06588__A1 _02752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05076_ _01567_ _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09953_ _00407_ io_in[4] u_cpu.rf_ram.memory\[54\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05260__A1 _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08329__A2 _03890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08904_ _04280_ _04309_ _04310_ _01077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09884_ _00338_ io_in[4] u_cpu.rf_ram.memory\[62\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07001__A2 _03071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08835_ _03811_ _03809_ _04266_ _04267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08766_ _02573_ u_cpu.rf_ram.memory\[2\]\[0\] _04217_ _04218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_57_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05978_ u_cpu.cpu.bufreg.c_r _02442_ _02443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_57_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06760__A1 _02744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07717_ _03349_ _03475_ _03478_ _00721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04929_ u_cpu.cpu.ctrl.o_ibus_adr\[4\] _01448_ _01449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_54_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08697_ _04178_ _01002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__08501__A2 _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07648_ _03355_ _03432_ _03438_ _00692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05315__A2 _01804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07579_ u_cpu.rf_ram.memory\[125\]\[7\] _03392_ _03400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09933__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09318_ u_cpu.rf_ram.memory\[111\]\[5\] _04536_ _04542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10590_ _01020_ io_in[4] u_cpu.rf_ram.memory\[109\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09249_ _04503_ _01229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10910__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06815__A2 _02727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08017__A1 u_arbiter.i_wb_cpu_dbus_dat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07240__A2 _03206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09517__A1 _04478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11073_ _11073_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_110_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10024_ _00470_ io_in[4] u_cpu.rf_ram.memory\[140\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[2\] u_arbiter.i_wb_cpu_ack io_in[3] u_arbiter.i_wb_cpu_dbus_sel\[0\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__05003__A1 _01445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08740__A2 _04199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05554__A2 _02041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10440__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10926_ _01354_ io_in[4] u_cpu.rf_ram.memory\[23\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06503__A1 _02742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05857__A3 _02338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10857_ _01286_ io_in[4] u_cpu.cpu.genblk3.csr.mstatus_mie vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08256__A1 _03763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08307__S _01436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10788_ _01217_ io_in[4] u_cpu.rf_ram.memory\[59\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10590__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08559__A2 _04094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07231__A2 _03196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06950_ u_cpu.rf_ram.memory\[57\]\[4\] _03041_ _03046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06070__B _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05901_ _02313_ _02383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09806__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06881_ u_cpu.rf_ram.memory\[60\]\[5\] _03002_ _03008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08620_ _04132_ _00971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05832_ _02306_ _02314_ u_cpu.cpu.immdec.imm24_20\[0\] _02316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_67_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06742__A1 _02744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08551_ _03545_ _04094_ _04097_ _00937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05763_ u_cpu.rf_ram.memory\[36\]\[7\] u_cpu.rf_ram.memory\[37\]\[7\] u_cpu.rf_ram.memory\[38\]\[7\]
+ u_cpu.rf_ram.memory\[39\]\[7\] _01619_ _01620_ _02248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09956__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07502_ _03355_ _03345_ _03356_ _00628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05414__B _01626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08482_ _04040_ _04043_ _04044_ _03940_ _04045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__07298__A2 _03235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05694_ _01601_ _02179_ _01605_ _02180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_35_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07433_ _03157_ _03315_ _03316_ _00599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10933__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08247__A1 _02332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07364_ u_cpu.rf_ram.memory\[135\]\[2\] _03275_ _03278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09103_ u_cpu.rf_ram.memory\[106\]\[0\] _04419_ _04420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06315_ u_cpu.rf_ram.memory\[44\]\[1\] _02673_ _02675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08798__A2 _04227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07295_ _03165_ _03235_ _03239_ _00538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09034_ _04284_ _04379_ _04381_ _01136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06246_ u_cpu.rf_ram.memory\[78\]\[5\] _02628_ _02634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06177_ _02589_ _02590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08460__B _03801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05128_ _01548_ _01620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07222__A2 _03196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10313__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05059_ u_cpu.rf_ram.memory\[8\]\[0\] u_cpu.rf_ram.memory\[9\]\[0\] u_cpu.rf_ram.memory\[10\]\[0\]
+ u_cpu.rf_ram.memory\[11\]\[0\] _01546_ _01550_ _01551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09936_ _00390_ io_in[4] u_cpu.rf_ram.memory\[57\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06981__A1 _02957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[9\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09867_ _00321_ io_in[4] u_cpu.rf_ram.memory\[29\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08722__A2 _01410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10463__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08818_ _03780_ _04249_ _04251_ _04024_ _04252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_73_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09798_ _00252_ io_in[4] u_cpu.rf_ram.memory\[74\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05092__S0 _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08749_ _02573_ u_cpu.rf_ram.memory\[3\]\[0\] _04208_ _04209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08486__A1 u_cpu.cpu.immdec.imm19_12_20\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07289__A2 _03235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10711_ _01140_ io_in[4] u_cpu.rf_ram.memory\[104\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05395__S1 _01580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10642_ _01071_ io_in[4] u_cpu.rf_ram.memory\[95\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08238__A1 _03825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08238__B2 _03801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08354__C _03797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08789__A2 _04227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10573_ _01003_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05147__S1 _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07461__A2 _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05994__B _02433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09829__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07213__A2 _03186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08410__A1 _03742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05775__A2 _02259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10806__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11056_ _11056_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_27_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09979__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10007_ _00453_ io_in[4] u_cpu.rf_ram.memory\[142\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06724__A1 _02744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05083__S0 _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10956__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05234__B _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08477__A1 _03747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10909_ _01338_ io_in[4] u_cpu.rf_ram.memory\[100\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05386__S1 _01557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08229__B2 _03757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06100_ _02540_ _02541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07080_ _02599_ u_cpu.rf_ram.memory\[15\]\[7\] _03109_ _03117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07452__A2 _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10336__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06031_ _02486_ _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08401__A1 _02765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07204__A2 _03186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07982_ _03551_ _03626_ _03632_ _00833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10486__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05195__I _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05310__S1 _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06963__A1 _02957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09721_ _00175_ io_in[4] u_cpu.rf_ram.memory\[50\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06933_ _02963_ _03031_ _03036_ _00379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08704__A2 _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09652_ _00106_ io_in[4] u_cpu.rf_ram.memory\[46\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06864_ _02965_ _02992_ _02998_ _00348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05518__A2 _02005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08439__C _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08603_ u_arbiter.i_wb_cpu_dbus_adr\[22\] u_arbiter.i_wb_cpu_dbus_adr\[21\] _04115_
+ _04124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05815_ u_cpu.rf_ram.memory\[132\]\[7\] u_cpu.rf_ram.memory\[133\]\[7\] u_cpu.rf_ram.memory\[134\]\[7\]
+ u_cpu.rf_ram.memory\[135\]\[7\] _01687_ _01688_ _02300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09583_ _00037_ io_in[4] u_cpu.rf_ram.memory\[21\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06795_ u_cpu.rf_ram.memory\[29\]\[1\] _02955_ _02958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08534_ u_cpu.rf_ram.memory\[32\]\[3\] _04084_ _04088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08468__A1 _03999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05746_ _01554_ _02230_ _02231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08465_ _03851_ _03896_ _04029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05677_ u_cpu.rf_ram.memory\[32\]\[6\] u_cpu.rf_ram.memory\[33\]\[6\] u_cpu.rf_ram.memory\[34\]\[6\]
+ u_cpu.rf_ram.memory\[35\]\[6\] _01623_ _01624_ _02163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_51_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07416_ u_cpu.rf_ram.memory\[132\]\[1\] _03305_ _03307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08396_ _02765_ u_arbiter.i_wb_cpu_rdt\[28\] _03967_ _03968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07347_ _03163_ _03265_ _03268_ _00561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05129__S1 _01620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07443__A2 _03315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07278_ u_cpu.rf_ram.memory\[138\]\[4\] _03225_ _03230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09017_ u_cpu.rf_ram.memory\[103\]\[2\] _04369_ _04372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06229_ _02517_ _02614_ _02622_ _00089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10829__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05757__A2 _02241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05301__S1 _01574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09919_ _00373_ io_in[4] u_cpu.rf_ram.memory\[5\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06706__A1 _02744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08171__A3 _03770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10209__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07131__A1 _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07682__A2 _02311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10359__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10625_ _01054_ io_in[4] u_cpu.rf_ram.memory\[97\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09651__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08631__A1 _02361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10556_ _00986_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07434__A2 _03315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10487_ _00920_ io_in[4] u_cpu.cpu.csr_imm vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05540__S1 _01549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09187__A2 _04459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05229__B _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08934__A2 _04322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06945__A1 _02957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05748__A2 _02232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11108_ io_oeb[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_96_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11039_ _11039_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_110_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05600_ u_cpu.rf_ram.memory\[96\]\[5\] u_cpu.rf_ram.memory\[97\]\[5\] u_cpu.rf_ram.memory\[98\]\[5\]
+ u_cpu.rf_ram.memory\[99\]\[5\] _01602_ _01579_ _02087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_40_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06580_ _02744_ _02834_ _02837_ _00225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_91_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05920__A2 _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09111__A2 _04419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05531_ u_cpu.rf_ram.memory\[84\]\[4\] u_cpu.rf_ram.memory\[85\]\[4\] u_cpu.rf_ram.memory\[86\]\[4\]
+ u_cpu.rf_ram.memory\[87\]\[4\] _01555_ _01652_ _02019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_127_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08250_ _03762_ _03790_ _03818_ _03842_ _03835_ _03843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_60_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05462_ _01399_ _01950_ _01951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08870__A1 _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07201_ u_cpu.rf_ram.memory\[71\]\[1\] _03186_ _03188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08181_ _03779_ _03780_ _03781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05393_ u_cpu.rf_ram.memory\[28\]\[3\] u_cpu.rf_ram.memory\[29\]\[3\] u_cpu.rf_ram.memory\[30\]\[3\]
+ u_cpu.rf_ram.memory\[31\]\[3\] _01572_ _01574_ _01882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07132_ u_cpu.rf_ram.memory\[140\]\[6\] _03139_ _03146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07425__A2 _03305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05436__A1 _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07063_ _02599_ u_cpu.rf_ram.memory\[9\]\[7\] _03100_ _03108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__05531__S1 _01652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06014_ u_cpu.rf_ram_if.genblk1.wtrig0_r u_cpu.rf_ram_if.wen1_r u_cpu.rf_ram_if.rtrig0
+ u_cpu.rf_ram_if.wen0_r _02471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09178__A2 _04459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07965_ u_cpu.rf_ram.memory\[115\]\[6\] _03616_ _03623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09704_ _00158_ io_in[4] u_cpu.rf_ram.memory\[48\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06916_ _02593_ u_cpu.rf_ram.memory\[5\]\[5\] _03021_ _03027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08689__A1 u_cpu.cpu.ctrl.o_ibus_adr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07896_ _02599_ u_cpu.rf_ram.memory\[8\]\[7\] _03577_ _03585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09350__A2 _04556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09635_ _00089_ io_in[4] u_cpu.rf_ram.memory\[80\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06847_ u_cpu.rf_ram.memory\[62\]\[6\] _02982_ _02989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07361__A1 _03157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05598__S1 _01549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06685__S _02894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09566_ _04686_ _01363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_70_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06778_ _02744_ _02944_ _02947_ _00313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10501__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08517_ _04016_ _04072_ _04075_ _04076_ _00924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_05729_ _02208_ _02210_ _02212_ _02214_ _01404_ _02215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_09497_ _04476_ _04644_ _04648_ _01332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07113__A1 _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09674__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08861__A1 _04280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07664__A2 _03442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08448_ _04015_ _04016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_141_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08379_ _03797_ _03948_ _03954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_104_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10410_ _00843_ io_in[4] u_cpu.rf_ram.memory\[33\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05770__S1 _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10651__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07416__A2 _03305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10341_ _00774_ io_in[4] u_cpu.rf_ram.memory\[118\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09169__A2 _04449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10272_ _00705_ io_in[4] u_cpu.cpu.mem_bytecnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08916__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06927__A1 _02957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09236__S _04496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10031__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09341__A2 _04546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05589__S1 _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08874__I _02506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10181__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08852__A1 _03551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07655__A2 _03442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05210__S0 _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05761__S1 _01616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10608_ _01037_ io_in[4] u_cpu.rf_ram.memory\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07407__A2 _03295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06466__I0 _02599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08080__A2 _03653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10539_ _00972_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06091__A1 _02502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08907__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09373__C _01375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06394__A2 _02718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07750_ _03343_ _03500_ _03501_ _00732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_04962_ u_cpu.cpu.ctrl.o_ibus_adr\[11\] u_cpu.cpu.ctrl.o_ibus_adr\[10\] _01475_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[22\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09332__A2 _04546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06701_ u_cpu.rf_ram.memory\[68\]\[0\] _02904_ _02905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10524__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07681_ _01428_ _03457_ _00706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04893_ u_cpu.cpu.immdec.imm19_12_20\[7\] _01368_ _01419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05406__C _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07343__A1 _03157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06146__A2 _02563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06632_ _02742_ _02864_ _02866_ _00248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09420_ _04468_ _04605_ _04606_ _01297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09697__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09351_ _04476_ _04556_ _04560_ _01274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06563_ _02746_ _02823_ _02827_ _00218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09096__A1 _04292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[37\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08143__I0 u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08302_ _03551_ _03879_ _03885_ _00900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05514_ _01995_ _01997_ _01999_ _02001_ _01628_ _02002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_21_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09282_ u_cpu.rf_ram.memory\[110\]\[5\] _04516_ _04522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10674__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07646__A2 _03432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06494_ _02769_ _02783_ _02786_ _02787_ _02788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_08233_ _03767_ _03778_ _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05445_ _01927_ _01929_ _01931_ _01933_ _01426_ _01934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_119_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05752__S1 _01548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08164_ _03761_ _03762_ _03763_ _03764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__09399__A2 _02706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05376_ _01684_ _01865_ _01418_ _01866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07115_ _02967_ _03129_ _03136_ _00461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08095_ _03711_ _03712_ _00866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07046_ u_cpu.rf_ram.memory\[52\]\[7\] _03091_ _03099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06209__I0 _02599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09020__A1 _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10054__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06385__A2 _02708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08997_ u_cpu.rf_ram.memory\[102\]\[1\] _04359_ _04361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07948_ _03553_ _03606_ _03613_ _00818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09323__A2 _04536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07879_ u_cpu.rf_ram.memory\[121\]\[7\] _03568_ _03576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06137__A2 _02561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09618_ _00072_ io_in[4] u_cpu.rf_ram.memory\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10890_ _01319_ io_in[4] u_cpu.rf_ram.memory\[24\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09549_ _04474_ _04674_ _04677_ _01355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_93_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07637__A2 _03432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[25\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05743__S1 _01557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10324_ _00757_ io_in[4] u_cpu.rf_ram.memory\[117\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10255_ _00688_ io_in[4] u_cpu.rf_ram.memory\[37\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09011__A1 _02602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09562__A2 _04683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10547__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10186_ _00632_ io_in[4] u_cpu.rf_ram.memory\[128\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06376__A2 _02708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09314__A2 _04536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06128__A2 _02551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07325__A1 _03157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10697__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07876__A2 _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05431__S0 _01619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09078__A1 _04292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07628__A2 _03422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06687__I0 _02584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06300__A2 _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05734__S1 _01668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05230_ _01714_ _01716_ _01718_ _01720_ _01607_ _01721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_128_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05161_ u_cpu.rf_ram.memory\[116\]\[0\] u_cpu.rf_ram.memory\[117\]\[0\] u_cpu.rf_ram.memory\[118\]\[0\]
+ u_cpu.rf_ram.memory\[119\]\[0\] _01623_ _01652_ _01653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_7_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04862__A2 _01377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10077__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07884__S _03577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06064__A1 _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05092_ u_cpu.rf_ram.memory\[28\]\[0\] u_cpu.rf_ram.memory\[29\]\[0\] u_cpu.rf_ram.memory\[30\]\[0\]
+ u_cpu.rf_ram.memory\[31\]\[0\] _01572_ _01574_ _01584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07800__A2 _03520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08920_ _03991_ _04318_ _01085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09002__A1 _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08851_ u_cpu.rf_ram.memory\[97\]\[5\] _04271_ _04277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09553__A2 _04674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06367__A2 _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07802_ _03529_ _03530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08782_ _02475_ _02660_ _04226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05994_ _01393_ _02454_ _02433_ u_cpu.cpu.o_wen0 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_85_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09305__A2 _04526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04945_ u_cpu.cpu.ctrl.o_ibus_adr\[8\] _01461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07733_ _02309_ _03487_ _03488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06119__A2 _02551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07867__A2 _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07664_ _03353_ _03442_ _03447_ _00699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_u_scanchain_local.scan_flop\[48\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04876_ _01400_ _01401_ _01402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05931__I _02411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05422__S0 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05878__A1 _01410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09403_ u_cpu.rf_ram.memory\[27\]\[1\] _04595_ _04597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06615_ u_cpu.rf_ram.memory\[77\]\[2\] _02854_ _02857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07595_ u_cpu.rf_ram.memory\[124\]\[6\] _03402_ _03409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09334_ u_cpu.rf_ram.memory\[87\]\[4\] _04546_ _04551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06546_ _02748_ _02812_ _02817_ _00211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07619__A2 _03422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08816__A1 _03743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09265_ _04480_ _04506_ _04512_ _01236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06477_ _02447_ _02365_ _02773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08292__A2 _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05725__S1 _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05428_ _01398_ _01916_ _01917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08216_ _03773_ _03767_ _03808_ _03813_ _03814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_14_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09196_ _02486_ _04472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_5_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09712__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08147_ _02765_ u_arbiter.i_wb_cpu_rdt\[8\] _03746_ _03747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05359_ _01667_ _01848_ _01849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08078_ u_arbiter.i_wb_cpu_rdt\[16\] _03669_ _03678_ u_arbiter.i_wb_cpu_dbus_dat\[16\]
+ _03702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_49_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07029_ _02969_ _03081_ _03089_ _00422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10040_ _00486_ io_in[4] u_cpu.rf_ram.memory\[72\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09862__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09544__A2 _04674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06203__S _02603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06358__A2 _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07307__A1 _03157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10942_ _01362_ io_in[4] u_cpu.rf_ram_if.rdata1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07858__A2 _03558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05869__A1 _02309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05413__S0 _01623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10873_ _01302_ io_in[4] u_cpu.rf_ram.memory\[26\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06530__A2 _02801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08807__A1 _03747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08807__B2 _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05997__B _02332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08283__A2 _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05716__S1 _01549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09232__A1 _04482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06046__A1 _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07794__A1 _03353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06597__A2 _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10307_ _00740_ io_in[4] u_cpu.rf_ram.memory\[35\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09535__A2 _04664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10238_ _00678_ io_in[4] u_cpu.rf_ram.memory\[123\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06349__A2 _02686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10169_ _00615_ io_in[4] u_cpu.rf_ram.memory\[12\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09299__A1 _04478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08346__I0 u_arbiter.i_wb_cpu_rdt\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07849__A2 _03558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05404__S0 _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06400_ u_cpu.rf_ram.memory\[48\]\[5\] _02718_ _02724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06521__A2 _02801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07380_ u_cpu.rf_ram.memory\[134\]\[1\] _03285_ _03287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06331_ _02526_ _02683_ _02684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_124_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09735__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09471__A1 _02577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05707__S1 _01652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09050_ _04280_ _04389_ _04390_ _01143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06262_ _02492_ _02641_ _02644_ _00100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08001_ u_cpu.rf_ram.memory\[33\]\[6\] _03636_ _03643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05213_ u_cpu.rf_ram.memory\[20\]\[1\] u_cpu.rf_ram.memory\[21\]\[1\] u_cpu.rf_ram.memory\[22\]\[1\]
+ u_cpu.rf_ram.memory\[23\]\[1\] _01572_ _01574_ _01704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_135_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10712__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06193_ _02523_ _02601_ _02602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09223__A1 u_cpu.rf_ram.memory\[59\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[0\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05144_ _01397_ _01636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09885__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06588__A2 _02834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05075_ _01423_ _01424_ _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09952_ _00406_ io_in[4] u_cpu.rf_ram.memory\[55\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10862__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09526__A2 _04664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08903_ u_cpu.rf_ram.memory\[96\]\[0\] _04309_ _04310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05260__A2 _01741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09883_ _00337_ io_in[4] u_cpu.rf_ram.memory\[62\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08834_ _03861_ _04265_ _03807_ _03851_ _04266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08765_ _02469_ _02577_ _04217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05977_ _02309_ _02437_ _02438_ _02442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_66_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06760__A2 _02934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07716_ u_cpu.rf_ram.memory\[90\]\[2\] _03475_ _03478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04928_ _01437_ u_cpu.cpu.ctrl.o_ibus_adr\[3\] u_cpu.cpu.ctrl.o_ibus_adr\[2\] _01448_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08696_ u_cpu.cpu.ctrl.o_ibus_adr\[18\] _04173_ _04175_ u_cpu.cpu.ctrl.o_ibus_adr\[19\]
+ _04178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_54_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07647_ u_cpu.rf_ram.memory\[37\]\[5\] _03432_ _03438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04859_ u_cpu.cpu.state.genblk1.misalign_trap_sync_r _01385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_80_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06512__A2 _02791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10242__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06693__S _02894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07578_ _03357_ _03392_ _03399_ _00661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09317_ _04478_ _04536_ _04541_ _01259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06529_ _02750_ _02801_ _02807_ _00204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09462__A1 _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06276__A1 _02482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05610__B _01654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09248_ _02596_ u_cpu.rf_ram.memory\[10\]\[6\] _04496_ _04503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10392__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08017__A2 _02774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09179_ u_cpu.rf_ram.memory\[69\]\[2\] _04459_ _04462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06028__A1 _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07076__I0 _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07776__A1 _03353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06579__A2 _02834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11072_ _11072_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__09517__A2 _04654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10023_ _00469_ io_in[4] u_cpu.rf_ram.memory\[140\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09608__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09244__S _04496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06751__A2 _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10925_ _01353_ io_in[4] u_cpu.rf_ram.memory\[23\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09758__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06503__A2 _02791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10856_ _01285_ io_in[4] u_cpu.cpu.genblk3.csr.mie_mtie vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05857__A4 _02339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10735__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08256__A2 _03785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09453__A1 _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10787_ _01216_ io_in[4] u_cpu.rf_ram.memory\[59\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04915__I _01436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06019__A1 _02469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10885__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09508__A2 _04654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10115__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08716__B1 _04175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06990__A2 _03061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05900_ _01374_ _02313_ _02382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06880_ _02963_ _03002_ _03007_ _00355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08192__A1 _03786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05831_ _02306_ _02312_ _02314_ _02315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_94_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06742__A2 _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10265__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05762_ _01397_ _02246_ _01416_ _02247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08550_ u_cpu.rf_ram.memory\[31\]\[2\] _04094_ _04097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07501_ u_cpu.rf_ram.memory\[22\]\[5\] _03345_ _03356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05693_ u_cpu.rf_ram.memory\[120\]\[6\] u_cpu.rf_ram.memory\[121\]\[6\] u_cpu.rf_ram.memory\[122\]\[6\]
+ u_cpu.rf_ram.memory\[123\]\[6\] _01646_ _01603_ _02179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08481_ _03747_ _03825_ _04026_ _03851_ _04044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_36_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08495__A2 _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07432_ u_cpu.rf_ram.memory\[131\]\[0\] _03315_ _03316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08247__A2 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07363_ _03161_ _03275_ _03277_ _00568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09444__A1 _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09102_ _04418_ _04419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06258__A1 _02482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05430__B _01648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06314_ _02482_ _02673_ _02674_ _00122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07294_ u_cpu.rf_ram.memory\[39\]\[3\] _03235_ _03239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09033_ u_cpu.rf_ram.memory\[104\]\[1\] _04379_ _04381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06245_ _02502_ _02628_ _02633_ _00094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06176_ u_cpu.rf_ram_if.wdata0_r\[4\] u_cpu.rf_ram_if.wdata1_r\[4\] _02478_ _02589_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_11_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07758__A1 _03353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05127_ _01544_ _01619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08032__I _03653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09935_ _00389_ io_in[4] u_cpu.rf_ram.memory\[57\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05058_ _01549_ _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06981__A2 _03061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__04992__A1 _01443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09866_ _00320_ io_in[4] u_cpu.rf_ram.memory\[29\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10608__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08183__A1 _03763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08817_ _03810_ _04250_ _03897_ _03873_ _04251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_85_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09797_ _00251_ io_in[4] u_cpu.rf_ram.memory\[74\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07930__A1 _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06733__A2 _02914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09900__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05092__S1 _01574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08748_ _02577_ _02682_ _04208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10758__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08679_ _04168_ _00994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__08486__A2 _04016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10710_ _01139_ io_in[4] u_cpu.rf_ram.memory\[104\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10641_ _01070_ io_in[4] u_cpu.rf_ram.memory\[95\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08238__A2 _03826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09435__A1 _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06249__A1 _02512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10572_ _01002_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07049__I0 _02573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08143__S _01435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10138__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08410__A2 _03786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06972__A2 _03051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10288__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11055_ _11055_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_122_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08877__I _02511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08174__A1 _03773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05607__S0 _01619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10006_ _00452_ io_in[4] u_cpu.rf_ram.memory\[142\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09580__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06724__A2 _02914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05083__S1 _01574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08477__A2 _03988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06488__A1 _02769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10908_ _01337_ io_in[4] u_cpu.rf_ram.memory\[100\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10839_ _01268_ io_in[4] u_cpu.rf_ram.memory\[87\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09426__A1 _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06030_ _02485_ _02486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06660__A1 _02752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08401__A2 u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07892__S _03577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06412__A1 _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07981_ u_cpu.rf_ram.memory\[116\]\[5\] _03626_ _03632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06963__A2 _03051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09923__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09720_ _00174_ io_in[4] u_cpu.rf_ram.memory\[50\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06932_ u_cpu.rf_ram.memory\[58\]\[4\] _03031_ _03036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__04974__A1 u_cpu.cpu.ctrl.o_ibus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08165__A1 _03757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09651_ _00105_ io_in[4] u_cpu.rf_ram.memory\[42\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06863_ u_cpu.rf_ram.memory\[61\]\[5\] _02992_ _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10900__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06715__A2 _02904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08602_ _04123_ _00962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05425__B _01626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05814_ _01570_ _02298_ _02299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09582_ _00036_ io_in[4] u_cpu.rf_ram.memory\[21\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06794_ _02486_ _02957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08533_ _03545_ _04084_ _04087_ _00929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05745_ u_cpu.rf_ram.memory\[28\]\[7\] u_cpu.rf_ram.memory\[29\]\[7\] u_cpu.rf_ram.memory\[30\]\[7\]
+ u_cpu.rf_ram.memory\[31\]\[7\] _01546_ _01550_ _02230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08468__A2 _03988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06479__A1 u_arbiter.i_wb_cpu_dbus_dat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08464_ _04024_ _04025_ _04027_ _04028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05676_ _01597_ _02161_ _02162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07415_ _03157_ _03305_ _03306_ _00591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09417__A1 _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08395_ _01437_ u_arbiter.i_wb_cpu_rdt\[12\] _03967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_11_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07346_ u_cpu.rf_ram.memory\[136\]\[2\] _03265_ _03268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07277_ _03165_ _03225_ _03229_ _00530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08640__A2 _04145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09016_ _04284_ _04369_ _04371_ _01128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05454__A2 _01938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06228_ u_cpu.rf_ram.memory\[80\]\[7\] _02614_ _02622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06159_ _02478_ _01386_ _02526_ _02575_ _02576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__10430__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06403__A1 _02512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06954__A2 _03041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09918_ _00372_ io_in[4] u_cpu.rf_ram.memory\[5\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__04965__A1 _01443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09849_ _00303_ io_in[4] u_cpu.rf_ram.memory\[65\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10580__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06706__A2 _02904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08951__I0 u_arbiter.i_wb_cpu_rdt\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05390__A1 _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07131__A2 _03139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06190__I0 _02599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09408__A1 _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10624_ _01053_ io_in[4] u_cpu.rf_ram.memory\[97\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06890__A1 _02953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10555_ _00985_ io_in[4] u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05445__A2 _01929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06642__A1 _02752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10486_ _00919_ io_in[4] u_cpu.cpu.immdec.imm19_12_20\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[32\] u_arbiter.i_wb_cpu_rdt\[29\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[26\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_6_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09946__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08395__A1 _01437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08601__S _04115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10923__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06945__A2 _03041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11107_ io_oeb[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_110_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08147__A1 _02765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11038_ _11038_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_65_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08698__A2 _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05245__B _01416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07370__A2 _03275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05381__A1 _01542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05530_ _01609_ _02017_ _02018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07122__A2 _03139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10303__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05461_ u_cpu.rf_ram.memory\[128\]\[3\] u_cpu.rf_ram.memory\[129\]\[3\] u_cpu.rf_ram.memory\[130\]\[3\]
+ u_cpu.rf_ram.memory\[131\]\[3\] _01687_ _01688_ _01950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_21_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08870__A2 _04282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07200_ _03157_ _03186_ _03187_ _00495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08180_ _03773_ _03755_ _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05392_ _01562_ _01880_ _01582_ _01881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07131_ _02965_ _03139_ _03145_ _00468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08083__B1 _03678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08622__A2 _02445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10453__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05436__A2 _01915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07062_ _03107_ _00437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06013_ u_cpu.cpu.immdec.imm11_7\[2\] _02457_ _02470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07189__A2 _03176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08386__A1 _03761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06936__A2 _03031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07964_ _03551_ _03616_ _03622_ _00825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09703_ _00157_ io_in[4] u_cpu.rf_ram.memory\[48\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06915_ _03026_ _00371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08689__A2 _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07895_ _03584_ _00794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09634_ _00088_ io_in[4] u_cpu.rf_ram.memory\[80\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_u_scanchain_local.scan_flop\[6\]_SI u_arbiter.i_wb_cpu_dbus_dat\[0\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06846_ _02965_ _02982_ _02988_ _00340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07361__A2 _03275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09565_ _02321_ u_cpu.rf_ram.rdata\[7\] u_cpu.rf_ram_if.rtrig0 _04686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__05372__A1 _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06777_ u_cpu.rf_ram.memory\[64\]\[2\] _02944_ _02947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08516_ u_cpu.cpu.immdec.imm19_12_20\[8\] _04016_ _04076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05728_ _01684_ _02213_ _01418_ _02214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09496_ u_cpu.rf_ram.memory\[98\]\[3\] _04644_ _04648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09819__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07113__A2 _03129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08447_ _02305_ _04014_ _02767_ _04015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05602__C _01628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05659_ u_cpu.rf_ram.memory\[24\]\[6\] u_cpu.rf_ram.memory\[25\]\[6\] u_cpu.rf_ram.memory\[26\]\[6\]
+ u_cpu.rf_ram.memory\[27\]\[6\] _01578_ _01580_ _02145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08861__A2 _04282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06872__A1 _02953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08378_ u_cpu.cpu.immdec.imm30_25\[1\] _03740_ _03949_ _03952_ _03953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_137_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09969__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07329_ _03163_ _03255_ _03258_ _00553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06624__A1 _02752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10340_ _00773_ io_in[4] u_cpu.rf_ram.memory\[118\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10946__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10271_ _00704_ io_in[4] u_cpu.cpu.state.o_cnt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08377__A1 _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06927__A2 _03031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04938__A1 _01431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08129__A1 _03545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07352__A2 _03265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10326__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05363__A1 _01667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07104__A2 _03129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08852__A2 _04271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10476__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05210__S1 _01557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10607_ _01036_ io_in[4] u_cpu.rf_ram.memory\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10538_ _00971_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06091__A2 _02530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10469_ _00902_ io_in[4] u_cpu.rf_ram.memory\[114\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08368__A1 _03831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07591__A2 _03402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04961_ u_cpu.cpu.ctrl.o_ibus_adr\[10\] _01471_ u_cpu.cpu.ctrl.o_ibus_adr\[11\] _01474_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_49_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06700_ _02903_ _02904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07680_ u_cpu.cpu.mem_bytecnt\[1\] _03456_ _03457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_04892_ _01417_ _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_65_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07343__A2 _03265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06631_ u_cpu.rf_ram.memory\[74\]\[1\] _02864_ _02866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05354__A1 _01609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09350_ u_cpu.rf_ram.memory\[88\]\[3\] _04556_ _04560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06562_ u_cpu.rf_ram.memory\[119\]\[3\] _02823_ _02827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10819__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09096__A2 _04409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08301_ u_cpu.rf_ram.memory\[114\]\[5\] _03879_ _03885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08143__I1 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05513_ _01601_ _02000_ _01626_ _02001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09281_ _04478_ _04516_ _04521_ _01243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06493_ _01680_ _02785_ _02787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__08843__A2 _04271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08232_ _03757_ _03759_ _03819_ _03827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06854__A1 _02953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05444_ _01553_ _01932_ _01654_ _01933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_140_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08163_ u_arbiter.i_wb_cpu_rdt\[2\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[2\]
+ _01435_ _03763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05375_ u_cpu.rf_ram.memory\[132\]\[2\] u_cpu.rf_ram.memory\[133\]\[2\] u_cpu.rf_ram.memory\[134\]\[2\]
+ u_cpu.rf_ram.memory\[135\]\[2\] _01687_ _01688_ _01865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07114_ u_cpu.rf_ram.memory\[141\]\[6\] _03129_ _03136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06606__A1 _02752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08094_ u_arbiter.i_wb_cpu_rdt\[22\] _03653_ _03654_ u_arbiter.i_wb_cpu_dbus_dat\[22\]
+ _03712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_106_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07045_ _02967_ _03091_ _03098_ _00429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06082__A2 _02530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09020__A2 _04369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08996_ _04280_ _04359_ _04360_ _01119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10349__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07947_ u_cpu.rf_ram.memory\[122\]\[6\] _03606_ _03613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05593__A1 _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07878_ _03553_ _03568_ _03575_ _00786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09641__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08531__A1 _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07334__A2 _03255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09617_ _00071_ io_in[4] u_cpu.rf_ram.memory\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06829_ u_cpu.rf_ram.memory\[63\]\[6\] _02972_ _02979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10499__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05896__A2 u_cpu.cpu.ctrl.i_iscomp vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09548_ u_cpu.rf_ram.memory\[23\]\[2\] _04674_ _04677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09087__A2 _04409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09791__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09479_ _04638_ _01324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_54_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10323_ _00756_ io_in[4] u_cpu.rf_ram.memory\[117\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_140_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10254_ _00687_ io_in[4] u_cpu.rf_ram.memory\[37\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09011__A2 _04197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10185_ _00631_ io_in[4] u_cpu.rf_ram.memory\[128\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07573__A2 _03392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05584__A1 _01609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07325__A2 _03255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05431__S1 _01620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09078__A2 _04399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07089__A1 _02959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08834__B _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06836__A1 _02953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07884__I0 _02581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05160_ _01547_ _01652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__04862__A3 _01387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05091_ _01562_ _01581_ _01582_ _01583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_144_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09002__A2 _04359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08850_ _03549_ _04271_ _04276_ _01057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09664__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07801_ _02524_ _02821_ _03529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08781_ _04225_ _01039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05575__A1 _01589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05993_ u_cpu.cpu.immdec.imm11_7\[4\] _02452_ _02453_ _02448_ _02454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07732_ _02334_ _02364_ _03487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_04944_ _01445_ _01459_ _01460_ u_arbiter.o_wb_cpu_adr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10641__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08513__A1 _01375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07316__A2 _03245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07663_ u_cpu.rf_ram.memory\[36\]\[4\] _03442_ _03447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05327__B2 _01816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04875_ u_cpu.cpu.immdec.imm24_20\[4\] _01388_ _01401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09402_ _04468_ _04595_ _04596_ _01289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06614_ _02742_ _02854_ _02856_ _00240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05422__S1 _01549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07594_ _03355_ _03402_ _03408_ _00668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09069__A2 _04399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09333_ _04476_ _04546_ _04550_ _01266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06545_ u_cpu.rf_ram.memory\[40\]\[4\] _02812_ _02817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10791__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08816__A2 _03826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09264_ u_cpu.rf_ram.memory\[85\]\[5\] _04506_ _04512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06476_ _01372_ _02332_ _02772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08215_ _03773_ _03810_ _03812_ _03813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_138_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05427_ u_cpu.rf_ram.memory\[124\]\[3\] u_cpu.rf_ram.memory\[125\]\[3\] u_cpu.rf_ram.memory\[126\]\[3\]
+ u_cpu.rf_ram.memory\[127\]\[3\] _01545_ _01642_ _01916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_53_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09195_ _04468_ _04470_ _04471_ _01207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10021__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08146_ _01436_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[8\] _03746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05358_ u_cpu.rf_ram.memory\[64\]\[2\] u_cpu.rf_ram.memory\[65\]\[2\] u_cpu.rf_ram.memory\[66\]\[2\]
+ u_cpu.rf_ram.memory\[67\]\[2\] _01571_ _01668_ _01848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_88_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08077_ u_arbiter.i_wb_cpu_dbus_dat\[17\] _03683_ _03701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05289_ _01773_ _01775_ _01777_ _01779_ _01404_ _01780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_07028_ u_cpu.rf_ram.memory\[53\]\[7\] _03081_ _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10171__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05653__I2 u_cpu.rf_ram.memory\[22\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07555__A2 _03382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05327__C _01628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08979_ u_cpu.rf_ram.memory\[101\]\[1\] _04349_ _04351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05566__A1 _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07307__A2 _03245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10941_ u_cpu.rf_ram_if.wtrig0 io_in[4] u_cpu.rf_ram_if.genblk1.wtrig0_r vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05413__S1 _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05869__A2 _02325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10872_ _01301_ io_in[4] u_cpu.rf_ram.memory\[26\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08807__A2 _03825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08654__B _01428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06818__A1 _02953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05177__S0 _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06294__A2 _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[21\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09232__A2 _04487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10514__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09687__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07794__A2 _03520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10306_ _00739_ io_in[4] u_cpu.rf_ram.memory\[92\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[36\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05518__B _01648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10237_ _00677_ io_in[4] u_cpu.rf_ram.memory\[123\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10664__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08743__A1 _03551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05557__A1 _01542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10168_ _00614_ io_in[4] u_cpu.rf_ram.memory\[130\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09299__A2 _04526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10099_ _00545_ io_in[4] u_cpu.rf_ram.memory\[137\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08346__I1 u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05309__A1 _01792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05404__S1 _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10044__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06330_ u_cpu.cpu.immdec.imm11_7\[2\] u_cpu.cpu.immdec.imm11_7\[3\] _02457_ _02683_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_128_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05168__S0 _01646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09471__A2 _02612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06285__A2 _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06261_ u_cpu.rf_ram.memory\[42\]\[2\] _02641_ _02644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08000_ _03551_ _03636_ _03642_ _00841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05212_ _01696_ _01698_ _01700_ _01702_ _01568_ _01703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_128_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10194__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[20\]_D u_arbiter.i_wb_cpu_rdt\[17\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_06192_ _02466_ _02520_ _02601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09223__A2 _04487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05143_ _01594_ _01634_ _01416_ _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07785__A2 _03520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08982__A1 _04286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05074_ _01562_ _01563_ _01565_ _01566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09951_ _00405_ io_in[4] u_cpu.rf_ram.memory\[55\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05796__A1 _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08902_ _04308_ _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05260__A3 _01750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09882_ _00336_ io_in[4] u_cpu.rf_ram.memory\[62\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07537__A2 _03372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[15\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08833_ _03773_ _03787_ _04265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05548__A1 _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08764_ _04216_ _01031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05976_ _01375_ _02356_ _02440_ _02441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_2708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07715_ _03347_ _03475_ _03477_ _00720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04927_ _01445_ _01446_ _01447_ u_arbiter.o_wb_cpu_adr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08695_ _04177_ _01001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_53_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05163__B _01654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07646_ _03353_ _03432_ _03437_ _00691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_04858_ u_cpu.cpu.genblk3.csr.o_new_irq _01384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_26_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07577_ u_cpu.rf_ram.memory\[125\]\[6\] _03392_ _03399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05720__A1 _02186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09316_ u_cpu.rf_ram.memory\[111\]\[4\] _04536_ _04541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06528_ u_cpu.rf_ram.memory\[17\]\[5\] _02801_ _02807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09462__A2 _04625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10537__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06276__A2 _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09247_ _04502_ _01228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_u_scanchain_local.scan_flop\[22\]_SI u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06459_ _02760_ _00181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08670__B1 _04157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_u_scanchain_local.scan_flop\[11\]_D u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09178_ _04284_ _04459_ _04461_ _01200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08129_ _03545_ _03731_ _03734_ _00878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10687__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07776__A2 _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05787__B2 _02271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11071_ _11071_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_27_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08725__A1 _02324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10022_ _00468_ io_in[4] u_cpu.rf_ram.memory\[140\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05539__A1 _01667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08489__B1 _03779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10067__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09150__A1 _04292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10924_ _00025_ io_in[4] u_cpu.rf_ram.regzero vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05398__S0 _01590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07700__A2 _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05711__A1 _01667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10855_ _01284_ io_in[4] u_cpu.cpu.genblk3.csr.mstatus_mpie vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05801__B _01654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10786_ _01215_ io_in[4] u_cpu.rf_ram.memory\[59\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08256__A3 _03809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09453__A2 _02810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06267__A2 _02641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xu_scanchain_local.scan_flop\[62\] u_scanchain_local.module_data_in\[61\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[24\] u_scanchain_local.clk u_scanchain_local.module_data_in\[62\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_12_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[9\]_D u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06019__A2 _02475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07767__A2 _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[38\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07519__A2 _03362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08192__A2 _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05830_ _01372_ u_cpu.cpu.decode.opcode\[1\] _02313_ _02314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_67_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05761_ u_cpu.rf_ram.memory\[44\]\[7\] u_cpu.rf_ram.memory\[45\]\[7\] u_cpu.rf_ram.memory\[46\]\[7\]
+ u_cpu.rf_ram.memory\[47\]\[7\] _01615_ _01616_ _02246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_82_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09702__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07500_ _02506_ _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08480_ _04030_ _04041_ _04042_ _04043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_39_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05692_ _01589_ _02177_ _02178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05389__S0 _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07431_ _03314_ _03315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05702__A1 _01398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07362_ u_cpu.rf_ram.memory\[135\]\[1\] _03275_ _03277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09852__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09444__A2 _04615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09101_ _02638_ _04197_ _04418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06313_ u_cpu.rf_ram.memory\[44\]\[0\] _02673_ _02674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06258__A2 _02641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07455__A1 _03163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05305__I1 u_cpu.rf_ram.memory\[29\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07293_ _03163_ _03235_ _03238_ _00537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09032_ _04280_ _04379_ _04380_ _01135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06244_ u_cpu.rf_ram.memory\[78\]\[4\] _02628_ _02633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06175_ _02588_ _00069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07758__A2 _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05126_ _01614_ _01617_ _01605_ _01618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__04841__I _01368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05769__A1 _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05057_ _01548_ _01549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09934_ _00388_ io_in[4] u_cpu.rf_ram.memory\[57\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09865_ _00319_ io_in[4] u_cpu.rf_ram.memory\[29\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08183__A2 _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09380__A1 _02311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08816_ _03743_ _03826_ _04250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06194__A1 _02577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09796_ _00250_ io_in[4] u_cpu.rf_ram.memory\[74\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07930__A2 _03596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08747_ _03555_ _04199_ _04207_ _01023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05959_ _01403_ _02418_ _02428_ _00012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05941__A1 _02321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09132__A1 _04292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08678_ u_cpu.cpu.ctrl.o_ibus_adr\[10\] _04155_ _04157_ u_cpu.cpu.ctrl.o_ibus_adr\[11\]
+ _04168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07629_ u_cpu.rf_ram.memory\[38\]\[5\] _03422_ _03428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10640_ _01069_ io_in[4] u_cpu.rf_ram.memory\[95\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06209__S _02603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09435__A2 _02695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06249__A2 _02628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10571_ _01001_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07997__A2 _03636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07749__A2 _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06421__A2 _02729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11054_ _11054_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_1_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09725__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08174__A2 _03755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10005_ _00451_ io_in[4] u_cpu.rf_ram.memory\[142\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05607__S1 _01620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07921__A2 _03596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[68\]_SI u_arbiter.o_wb_cpu_adr\[30\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10702__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05932__A1 _02321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09875__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08826__C _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10907_ _01336_ io_in[4] u_cpu.rf_ram.memory\[98\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06488__A2 _02783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10838_ _01267_ io_in[4] u_cpu.rf_ram.memory\[87\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10852__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05791__S0 _01646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09426__A2 _04605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07437__A1 _03163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05250__C _01628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10769_ _01198_ io_in[4] u_cpu.rf_ram.memory\[108\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05999__A1 _01386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06660__A2 _02874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08937__A1 _04292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06412__A2 _02729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07980_ _03549_ _03626_ _03631_ _00832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_141_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10232__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06931_ _02961_ _03031_ _03035_ _00378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08165__A2 _03759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09650_ _00104_ io_in[4] u_cpu.rf_ram.memory\[42\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06862_ _02963_ _02992_ _02997_ _00347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08601_ u_arbiter.i_wb_cpu_dbus_adr\[21\] u_arbiter.i_wb_cpu_dbus_adr\[20\] _04115_
+ _04123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05813_ u_cpu.rf_ram.memory\[128\]\[7\] u_cpu.rf_ram.memory\[129\]\[7\] u_cpu.rf_ram.memory\[130\]\[7\]
+ u_cpu.rf_ram.memory\[131\]\[7\] _01572_ _01574_ _02298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10382__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09581_ _00035_ io_in[4] u_cpu.rf_ram.memory\[21\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06793_ _02953_ _02955_ _02956_ _00319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09114__A1 _04292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08532_ u_cpu.rf_ram.memory\[32\]\[2\] _04084_ _04087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05744_ _01562_ _02228_ _01582_ _02229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_36_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06479__A2 u_arbiter.i_wb_cpu_dbus_dat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08463_ _03825_ _03776_ _04026_ _04027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__07676__A1 _01428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05675_ u_cpu.rf_ram.memory\[36\]\[6\] u_cpu.rf_ram.memory\[37\]\[6\] u_cpu.rf_ram.memory\[38\]\[6\]
+ u_cpu.rf_ram.memory\[39\]\[6\] _01619_ _01620_ _02161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_51_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07414_ u_cpu.rf_ram.memory\[132\]\[0\] _03305_ _03306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08394_ _03965_ _03966_ _00911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09417__A2 _02638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07345_ _03161_ _03265_ _03267_ _00560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07979__A2 _03626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07276_ u_cpu.rf_ram.memory\[138\]\[3\] _03225_ _03229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05534__S0 _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09015_ u_cpu.rf_ram.memory\[103\]\[1\] _04369_ _04371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08471__C _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06227_ _02512_ _02614_ _02621_ _00088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06651__A2 _02874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06158_ _02470_ _02574_ _02575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09748__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05109_ _01540_ _01601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_104_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06403__A2 _02718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06089_ _02497_ _02530_ _02534_ _00037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05611__B1 _02095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09917_ _00371_ io_in[4] u_cpu.rf_ram.memory\[5\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10725__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09353__A1 _04478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05616__B _01648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09848_ _00302_ io_in[4] u_cpu.rf_ram.memory\[66\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09898__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09779_ _00233_ io_in[4] u_cpu.rf_ram.memory\[139\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10875__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05390__A2 _01878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09408__A2 _04595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10105__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10623_ _01052_ io_in[4] u_cpu.cpu.immdec.imm11_7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07419__A1 _03163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06890__A2 _03012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10554_ _00984_ io_in[4] u_arbiter.i_wb_cpu_ibus_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05525__S0 _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06642__A2 _02864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10485_ _00918_ io_in[4] u_cpu.cpu.immdec.imm19_12_20\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10255__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08919__A1 u_cpu.cpu.bufreg.i_sh_signed vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08395__A2 u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[25\] u_arbiter.i_wb_cpu_rdt\[22\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[19\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_111_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05602__B1 _02086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11106_ io_oeb[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_1_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08147__A2 u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11037_ _11037_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_110_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05381__A2 _01869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07658__A1 _03347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05460_ _01684_ _01948_ _01582_ _01949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06330__A1 u_cpu.cpu.immdec.imm11_7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06881__A2 _03002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05391_ u_cpu.rf_ram.memory\[16\]\[3\] u_cpu.rf_ram.memory\[17\]\[3\] u_cpu.rf_ram.memory\[18\]\[3\]
+ u_cpu.rf_ram.memory\[19\]\[3\] _01578_ _01580_ _01880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07130_ u_cpu.rf_ram.memory\[140\]\[5\] _03139_ _03145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08083__A1 u_arbiter.i_wb_cpu_rdt\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07061_ _02596_ u_cpu.rf_ram.memory\[9\]\[6\] _03100_ _03107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__05436__A3 _01924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06633__A2 _02864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06012_ _02464_ _02468_ _02469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10748__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08386__A2 _03860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06397__A1 _02497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07963_ u_cpu.rf_ram.memory\[115\]\[5\] _03616_ _03622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__04947__A2 _01462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08138__A2 _03731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09335__A1 _04478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06914_ _02590_ u_cpu.rf_ram.memory\[5\]\[4\] _03021_ _03026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09702_ _00156_ io_in[4] u_cpu.rf_ram.memory\[48\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07894_ _02596_ u_cpu.rf_ram.memory\[8\]\[6\] _03577_ _03584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10898__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09633_ _00087_ io_in[4] u_cpu.rf_ram.memory\[80\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06845_ u_cpu.rf_ram.memory\[62\]\[5\] _02982_ _02988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09564_ _04685_ _01362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06776_ _02742_ _02944_ _02946_ _00312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07143__S _03148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10128__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08515_ _01374_ _02392_ _04074_ _04075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_130_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05727_ u_cpu.rf_ram.memory\[132\]\[6\] u_cpu.rf_ram.memory\[133\]\[6\] u_cpu.rf_ram.memory\[134\]\[6\]
+ u_cpu.rf_ram.memory\[135\]\[6\] _01687_ _01688_ _02213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09495_ _04474_ _04644_ _04647_ _01331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08310__A2 _03788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08446_ _02317_ _02391_ _04013_ _04014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_51_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05658_ _01570_ _02143_ _02144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08377_ _03816_ _03950_ _03951_ _03952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06872__A2 _03002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05589_ u_cpu.rf_ram.memory\[32\]\[5\] u_cpu.rf_ram.memory\[33\]\[5\] u_cpu.rf_ram.memory\[34\]\[5\]
+ u_cpu.rf_ram.memory\[35\]\[5\] _01623_ _01624_ _02076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10278__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04883__A1 _01370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07328_ u_cpu.rf_ram.memory\[49\]\[2\] _03255_ _03258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08074__A1 u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06624__A2 _02854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07259_ _03219_ _00522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10270_ _00703_ io_in[4] u_cpu.cpu.state.stage_two_req vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06388__A1 _02612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08129__A2 _03731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05060__A1 _01542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05346__B _01654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06021__I u_cpu.rf_ram_if.genblk1.wtrig0_r vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05363__A2 _01852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07053__S _03100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05860__I u_cpu.cpu.decode.op21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08301__A2 _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09913__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06863__A2 _02992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10606_ _01035_ io_in[4] u_cpu.rf_ram.memory\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07812__A1 _03353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10537_ _00970_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06615__A2 _02854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10468_ _00901_ io_in[4] u_cpu.rf_ram.memory\[114\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09565__A1 _02321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10399_ _00832_ io_in[4] u_cpu.rf_ram.memory\[116\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06379__A1 _02497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07040__A2 _03091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09317__A1 _04478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04960_ _01469_ _01473_ u_arbiter.o_wb_cpu_adr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04891_ _01416_ _01417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08540__A2 _04084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06630_ _02738_ _02864_ _02865_ _00247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_92_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06561_ _02744_ _02823_ _02826_ _00217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_64_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08300_ _03549_ _03879_ _03884_ _00899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05512_ u_cpu.rf_ram.memory\[96\]\[4\] u_cpu.rf_ram.memory\[97\]\[4\] u_cpu.rf_ram.memory\[98\]\[4\]
+ u_cpu.rf_ram.memory\[99\]\[4\] _01602_ _01579_ _02000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09280_ u_cpu.rf_ram.memory\[110\]\[4\] _04516_ _04521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10420__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06303__A1 _02502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06492_ _01680_ _02785_ _02786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08231_ _03767_ _03778_ _03826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09593__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05443_ u_cpu.rf_ram.memory\[84\]\[3\] u_cpu.rf_ram.memory\[85\]\[3\] u_cpu.rf_ram.memory\[86\]\[3\]
+ u_cpu.rf_ram.memory\[87\]\[3\] _01555_ _01652_ _01932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06854__A2 _02992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04865__A1 _01390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08162_ u_arbiter.i_wb_cpu_rdt\[4\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[4\]
+ _01435_ _03762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05374_ _01399_ _01863_ _01864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10570__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07113_ _02965_ _03129_ _03135_ _00460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08093_ u_arbiter.i_wb_cpu_dbus_dat\[23\] _03683_ _03711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06606__A2 _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07044_ u_cpu.rf_ram.memory\[52\]\[6\] _03091_ _03098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05290__A1 _01771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08995_ u_cpu.rf_ram.memory\[102\]\[0\] _04359_ _04360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07946_ _03551_ _03606_ _03612_ _00817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05593__A2 _02051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06790__A1 _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07877_ u_cpu.rf_ram.memory\[121\]\[6\] _03568_ _03575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08477__B _03801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08531__A2 _04084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09616_ _00070_ io_in[4] u_cpu.rf_ram.memory\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06828_ _02965_ _02972_ _02978_ _00332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06542__A1 _02744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09547_ _04472_ _04674_ _04676_ _01354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06759_ u_cpu.rf_ram.memory\[65\]\[2\] _02934_ _02937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09936__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07098__A2 _03119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09478_ _02587_ u_cpu.rf_ram.memory\[0\]\[3\] _04634_ _04638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_24_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08429_ _01436_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[7\] _03998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__06845__A2 _02982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10913__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04856__A1 u_cpu.cpu.decode.op21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10322_ _00755_ io_in[4] u_cpu.rf_ram.memory\[34\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07270__A2 _03225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09547__A1 _04472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10253_ _00686_ io_in[4] u_cpu.rf_ram.memory\[38\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07022__A2 _03081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10184_ _00630_ io_in[4] u_cpu.rf_ram.memory\[22\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05033__A1 _01445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05584__A2 _02070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06908__I0 _02581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10443__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06533__A1 _02754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05523__C _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08286__A1 _03796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07089__A2 _03119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08607__S _04115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10593__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08834__C _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06836__A2 _02982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08038__A1 _02774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05090_ _01565_ _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09809__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08210__A1 _03752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07800_ _03359_ _03520_ _03528_ _00755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08780_ _02599_ u_cpu.rf_ram.memory\[2\]\[7\] _04217_ _04225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05992_ _02306_ _02313_ _02382_ _01373_ _02453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__05575__A2 _02061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07731_ u_cpu.cpu.ctrl.i_jump _03458_ _03486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04943_ u_arbiter.i_wb_cpu_dbus_adr\[7\] _01457_ _01460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09959__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08513__A2 u_cpu.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07662_ _03351_ _03442_ _03446_ _00698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_77_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04874_ u_cpu.cpu.immdec.imm19_12_20\[8\] _01368_ _01400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09401_ u_cpu.rf_ram.memory\[27\]\[0\] _04595_ _04596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06613_ u_cpu.rf_ram.memory\[77\]\[1\] _02854_ _02856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07593_ u_cpu.rf_ram.memory\[124\]\[5\] _03402_ _03408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10936__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06544_ _02746_ _02812_ _02816_ _00210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09332_ u_cpu.rf_ram.memory\[87\]\[3\] _04546_ _04550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09263_ _04478_ _04506_ _04511_ _01235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06475_ u_arbiter.i_wb_cpu_dbus_dat\[6\] _02770_ _02771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06827__A2 _02972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08214_ _02768_ _03811_ _03812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05426_ _01908_ _01910_ _01912_ _01914_ _01628_ _01915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_18_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08029__A1 u_arbiter.i_wb_cpu_rdt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09194_ u_cpu.rf_ram.memory\[84\]\[0\] _04470_ _04471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08145_ _03741_ _03742_ _03743_ _03744_ _03745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_05357_ _01840_ _01842_ _01844_ _01846_ _01426_ _01847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_135_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08076_ _03699_ _03700_ _00859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05288_ _01684_ _01778_ _01418_ _01779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10316__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09529__A1 _04472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07027_ _02967_ _03081_ _03088_ _00421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08201__A1 _02765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07004__A2 _03071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10466__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08978_ _04280_ _04349_ _04350_ _01111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07929_ u_cpu.rf_ram.memory\[112\]\[6\] _03596_ _03603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08504__A2 _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10940_ u_cpu.cpu.o_wdata0 io_in[4] u_cpu.rf_ram_if.wdata0_r\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06515__A1 _02754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10871_ _01300_ io_in[4] u_cpu.rf_ram.memory\[26\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08268__A1 _03773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06818__A2 _02972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05177__S1 _01668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08162__S _01435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07243__A2 _03206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05254__A1 _01645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10305_ _00738_ io_in[4] u_cpu.rf_ram.memory\[92\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08991__A2 _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10809__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10236_ _00676_ io_in[4] u_cpu.rf_ram.memory\[123\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09240__I0 _02584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08743__A2 _04199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10167_ _00613_ io_in[4] u_cpu.rf_ram.memory\[130\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05557__A2 _02043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10098_ _00544_ io_in[4] u_cpu.rf_ram.memory\[137\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08259__A1 _03754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05168__S1 _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06260_ _02487_ _02641_ _02643_ _00099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10339__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05211_ _01562_ _01701_ _01565_ _01702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05493__A1 _01601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06191_ _02600_ _00073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05142_ u_cpu.rf_ram.memory\[104\]\[0\] u_cpu.rf_ram.memory\[105\]\[0\] u_cpu.rf_ram.memory\[106\]\[0\]
+ u_cpu.rf_ram.memory\[107\]\[0\] _01615_ _01616_ _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09631__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08431__A1 _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05245__A1 _01594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08982__A2 _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05073_ _01564_ _01565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09950_ _00404_ io_in[4] u_cpu.rf_ram.memory\[55\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10489__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05796__A2 _02280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06993__A1 _02969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08901_ _02612_ _04197_ _04308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09881_ _00335_ io_in[4] u_cpu.rf_ram.memory\[62\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09781__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08734__A2 _04199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08832_ _04264_ _01051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05975_ u_cpu.cpu.decode.opcode\[1\] _02313_ _02440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08763_ _02599_ u_cpu.rf_ram.memory\[3\]\[7\] _04208_ _04216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_73_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07714_ u_cpu.rf_ram.memory\[90\]\[1\] _03475_ _03477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05444__B _01654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04926_ u_arbiter.i_wb_cpu_dbus_adr\[3\] _01443_ _01447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08694_ u_cpu.cpu.ctrl.o_ibus_adr\[17\] _04173_ _04175_ u_cpu.cpu.ctrl.o_ibus_adr\[18\]
+ _04177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_26_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07645_ u_cpu.rf_ram.memory\[37\]\[4\] _03432_ _03437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04857_ _01369_ _01370_ u_cpu.cpu.decode.op21 u_cpu.cpu.bne_or_bge _01383_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_53_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07576_ _03355_ _03392_ _03398_ _00660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07151__S _03148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09315_ _04476_ _04536_ _04540_ _01258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06527_ _02748_ _02801_ _02806_ _00203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06458_ _02587_ u_cpu.rf_ram.memory\[4\]\[3\] _02756_ _02760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09246_ _02593_ u_cpu.rf_ram.memory\[10\]\[5\] _04496_ _04502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_142_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05484__A1 _01542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05409_ u_cpu.rf_ram.memory\[44\]\[3\] u_cpu.rf_ram.memory\[45\]\[3\] u_cpu.rf_ram.memory\[46\]\[3\]
+ u_cpu.rf_ram.memory\[47\]\[3\] _01615_ _01616_ _01898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_108_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09177_ u_cpu.rf_ram.memory\[69\]\[1\] _04459_ _04461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06389_ _02717_ _02718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08128_ u_cpu.rf_ram.memory\[113\]\[2\] _03731_ _03734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07225__A2 _03196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05236__A1 _01589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08059_ _03688_ _03689_ _00853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11070_ _11070_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05338__C _01628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10021_ _00467_ io_in[4] u_cpu.rf_ram.memory\[140\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08725__A2 _02356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05539__A2 _02026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08489__A1 _03743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09150__A2 _04439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10923_ _01352_ io_in[4] u_cpu.rf_ram.memory\[89\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05398__S1 _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10854_ _01283_ io_in[4] u_cpu.cpu.genblk3.csr.mcause31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05711__A2 _02196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07061__S _03100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10785_ _01214_ io_in[4] u_cpu.rf_ram.memory\[84\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09654__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07464__A2 _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05475__A1 _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[55\] u_scanchain_local.module_data_in\[54\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[17\] u_scanchain_local.clk u_scanchain_local.module_data_in\[55\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__10631__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05227__A1 _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06975__A1 _02969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10781__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08716__A2 _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10219_ _00665_ io_in[4] u_cpu.rf_ram.memory\[124\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10011__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05264__B _01648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05760_ _01609_ _02244_ _02245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05950__A2 _01403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09141__A2 _04439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05691_ u_cpu.rf_ram.memory\[124\]\[6\] u_cpu.rf_ram.memory\[125\]\[6\] u_cpu.rf_ram.memory\[126\]\[6\]
+ u_cpu.rf_ram.memory\[127\]\[6\] _01545_ _01642_ _02177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_36_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05389__S1 _01574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07430_ _02682_ _02832_ _03314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10161__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07361_ _03157_ _03275_ _03276_ _00567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06312_ _02672_ _02673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09100_ _04296_ _04409_ _04417_ _01166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07455__A2 _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07292_ u_cpu.rf_ram.memory\[39\]\[2\] _03235_ _03238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09031_ u_cpu.rf_ram.memory\[104\]\[0\] _04379_ _04380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05466__A1 _01945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06243_ _02497_ _02628_ _02632_ _00093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07207__A2 _03186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08404__A1 _02305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06174_ _02587_ u_cpu.rf_ram.memory\[1\]\[3\] _02578_ _02588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05218__A1 _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05125_ u_cpu.rf_ram.memory\[44\]\[0\] u_cpu.rf_ram.memory\[45\]\[0\] u_cpu.rf_ram.memory\[46\]\[0\]
+ u_cpu.rf_ram.memory\[47\]\[0\] _01615_ _01616_ _01617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_102_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05769__A2 _02225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05056_ _01547_ _01548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09933_ _00387_ io_in[4] u_cpu.rf_ram.memory\[57\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09864_ _00318_ io_in[4] u_cpu.rf_ram.memory\[64\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08469__C _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08815_ _03973_ _03769_ _03809_ _03757_ _04248_ _04249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__09380__A2 _02344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09795_ _00249_ io_in[4] u_cpu.rf_ram.memory\[74\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06194__A2 _02602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07391__A1 _03171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08746_ u_cpu.rf_ram.memory\[109\]\[7\] _04199_ _04207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[20\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05958_ u_cpu.rf_ram_if.rdata0\[5\] _01403_ _02428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09132__A2 _04429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04909_ _01432_ u_arbiter.o_wb_cpu_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10504__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08677_ _04167_ _00993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_05889_ _02366_ _02370_ _02371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_57_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07628_ _03353_ _03422_ _03427_ _00683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09677__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07694__A2 _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[35\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07559_ u_cpu.rf_ram.memory\[126\]\[6\] _03382_ _03389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05621__C _01426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10654__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10570_ _01000_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07446__A2 _03315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08643__A1 _03545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09229_ u_cpu.rf_ram.memory\[59\]\[5\] _04487_ _04493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05209__A1 _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06957__A1 _02969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11053_ _11053_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_67_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10034__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05068__S0 _01546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10004_ _00450_ io_in[4] u_cpu.rf_ram.memory\[142\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[0\] io_in[2] io_in[3] u_arbiter.o_wb_cpu_cyc u_scanchain_local.clk
+ u_cpu.cpu.genblk3.csr.i_mtip vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_67_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09123__A2 _04429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10184__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10906_ _01335_ io_in[4] u_cpu.rf_ram.memory\[98\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05812__B _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08882__A1 _04296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05696__A1 _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10837_ _01266_ io_in[4] u_cpu.rf_ram.memory\[87\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05791__S1 _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07437__A2 _03315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10768_ _01197_ io_in[4] u_cpu.rf_ram.memory\[108\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08615__S _04115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10699_ _01128_ io_in[4] u_cpu.rf_ram.memory\[103\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05999__A2 _01394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08398__B1 _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08937__A2 _04322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05620__A1 _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06930_ u_cpu.rf_ram.memory\[58\]\[3\] _03031_ _03035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05059__S0 _01546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10527__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06861_ u_cpu.rf_ram.memory\[61\]\[4\] _02992_ _02997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[12\]_SI u_arbiter.i_wb_cpu_dbus_dat\[6\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07373__A1 _03171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08600_ _04122_ _00961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05812_ _01684_ _02296_ _01582_ _02297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06792_ u_cpu.rf_ram.memory\[29\]\[0\] _02955_ _02956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09580_ _00034_ io_in[4] u_cpu.rf_ram.memory\[21\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09114__A2 _04419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08531_ _03543_ _04084_ _04086_ _00928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05743_ u_cpu.rf_ram.memory\[16\]\[7\] u_cpu.rf_ram.memory\[17\]\[7\] u_cpu.rf_ram.memory\[18\]\[7\]
+ u_cpu.rf_ram.memory\[19\]\[7\] _01556_ _01557_ _02228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07125__A1 _02959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10677__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05674_ _01397_ _02159_ _01416_ _02160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08462_ _03751_ _03765_ _03768_ _04026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_35_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08873__A1 _04290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06479__A3 u_arbiter.i_wb_cpu_dbus_dat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05687__A1 _01636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05231__S0 _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07413_ _03304_ _03305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08393_ u_cpu.cpu.immdec.imm30_25\[2\] _03954_ _03956_ u_cpu.cpu.immdec.imm30_25\[3\]
+ _03963_ _03816_ _03966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_51_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07344_ u_cpu.rf_ram.memory\[136\]\[1\] _03265_ _03267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08625__A1 _01372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07428__A2 _03305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07275_ _03163_ _03225_ _03228_ _00529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05534__S1 _01668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09014_ _04280_ _04369_ _04370_ _01127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06226_ u_cpu.rf_ram.memory\[80\]\[6\] _02614_ _02621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08389__B1 _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05169__B _01648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06157_ u_cpu.cpu.immdec.imm11_7\[3\] _02457_ _02574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08928__A2 _04322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10057__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09050__A1 _04280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06939__A1 _02969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05298__S0 _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05108_ _01597_ _01599_ _01600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06088_ u_cpu.rf_ram.memory\[21\]\[3\] _02530_ _02534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05611__A1 _02091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09916_ _00370_ io_in[4] u_cpu.rf_ram.memory\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05039_ u_cpu.cpu.ctrl.o_ibus_adr\[30\] _01532_ _01533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_99_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09353__A2 _04556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09847_ _00301_ io_in[4] u_cpu.rf_ram.memory\[66\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09778_ _00232_ io_in[4] u_cpu.rf_ram.memory\[139\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05914__A2 u_cpu.cpu.mem_bytecnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09105__A2 _04419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05470__S0 _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08729_ u_cpu.cpu.immdec.imm11_7\[2\] _02473_ _02574_ _04197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05632__B _01402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08864__A1 _04284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07667__A2 _03442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[28\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07911__I0 _02596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05678__A1 _01645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05222__S0 _01590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10622_ _01051_ io_in[4] u_cpu.cpu.immdec.imm11_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07419__A2 _03305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10553_ _00023_ io_in[4] u_cpu.cpu.ctrl.pc_plus_4_cy_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05525__S1 _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10484_ _00917_ io_in[4] u_cpu.cpu.immdec.imm19_12_20\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08919__A2 _03798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11105_ io_oeb[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[18\] u_arbiter.i_wb_cpu_rdt\[15\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[12\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_89_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09344__A2 _04556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09842__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11036_ _11036_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__07355__A1 _03171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05461__S0 _01687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07741__C _01374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07107__A1 _02959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08155__I0 u_arbiter.i_wb_cpu_rdt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09992__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07658__A2 _03442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05213__S0 _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05669__A1 _01601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06330__A2 u_cpu.cpu.immdec.imm11_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05390_ _01570_ _01878_ _01879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08083__A2 _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07060_ _03106_ _00436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_12_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06011_ _01591_ _02467_ _02468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09032__A1 _04280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07594__A1 _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06397__A2 _02718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07962_ _03549_ _03616_ _03621_ _00824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05717__B _01648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09701_ _00155_ io_in[4] u_cpu.rf_ram.memory\[48\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09335__A2 _04546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06913_ _03025_ _00370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07893_ _03583_ _00793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06149__A2 _02563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09632_ _00086_ io_in[4] u_cpu.rf_ram.memory\[80\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06844_ _02963_ _02982_ _02987_ _00339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05452__S0 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09563_ _02321_ _02320_ u_cpu.rf_ram.rdata\[7\] _04685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_06775_ u_cpu.rf_ram.memory\[64\]\[1\] _02944_ _02946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08514_ _03797_ _04073_ _04074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__04847__I _01372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05726_ _01399_ _02211_ _02212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_64_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09494_ u_cpu.rf_ram.memory\[98\]\[2\] _04644_ _04647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08846__A1 _03545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07649__A2 _03432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05204__S0 _01546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08445_ _01373_ u_cpu.cpu.decode.opcode\[1\] _04013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05657_ u_cpu.rf_ram.memory\[28\]\[6\] u_cpu.rf_ram.memory\[29\]\[6\] u_cpu.rf_ram.memory\[30\]\[6\]
+ u_cpu.rf_ram.memory\[31\]\[6\] _01546_ _01574_ _02143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06321__A2 _02673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05588_ _01597_ _02074_ _02075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08376_ _01437_ u_arbiter.i_wb_cpu_rdt\[9\] _03951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08482__C _03940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09715__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04883__A2 u_cpu.cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07327_ _03161_ _03255_ _03257_ _00552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08074__A2 _03683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06085__A1 _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07258_ _02587_ u_cpu.rf_ram.memory\[14\]\[3\] _03215_ _03219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__05832__A1 _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06209_ _02599_ u_cpu.rf_ram.memory\[7\]\[7\] _02603_ _02611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07189_ u_cpu.rf_ram.memory\[73\]\[4\] _03176_ _03181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09865__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06388__A2 _02684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10842__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09326__A2 _04546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05060__A2 _01551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05691__S0 _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07337__A1 _03171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05443__S0 _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06560__A2 _02823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08837__A1 u_cpu.cpu.immdec.imm30_25\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10222__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10605_ _01034_ io_in[4] u_cpu.rf_ram.memory\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__04874__A2 _01368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10536_ _00969_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07812__A2 _03530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10372__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09014__A1 _04280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10467_ _00900_ io_in[4] u_cpu.rf_ram.memory\[114\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07576__A1 _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10398_ _00831_ io_in[4] u_cpu.rf_ram.memory\[116\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06379__A2 _02708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05537__B _01565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09317__A2 _04536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05682__S0 _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11019_ _11019_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_93_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04890_ _01415_ _01416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07879__A2 _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06000__A1 u_cpu.rf_ram_if.genblk1.wtrig0_r vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06551__A2 _02812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06560_ u_cpu.rf_ram.memory\[119\]\[2\] _02823_ _02826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08828__A1 _03801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05511_ _01636_ _01998_ _01999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06491_ _02465_ _02784_ _02785_ _00188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__09738__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06303__A2 _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05442_ _01609_ _01930_ _01931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08230_ _03754_ _03755_ _03825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10715__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04865__A2 u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08161_ _01435_ _03668_ _03760_ _03761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05373_ u_cpu.rf_ram.memory\[128\]\[2\] u_cpu.rf_ram.memory\[129\]\[2\] u_cpu.rf_ram.memory\[130\]\[2\]
+ u_cpu.rf_ram.memory\[131\]\[2\] _01687_ _01688_ _01863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07112_ u_cpu.rf_ram.memory\[141\]\[5\] _03129_ _03135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08092_ _03710_ _00865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__09888__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07803__A2 _03530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07043_ _02965_ _03091_ _03097_ _00428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05814__A1 _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10865__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09556__A2 _04674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05290__A2 _01780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08994_ _04358_ _04359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09308__A2 _04536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05673__S0 _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07945_ u_cpu.rf_ram.memory\[122\]\[5\] _03606_ _03612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07319__A1 _03171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05593__A3 _02060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06790__A2 _02660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07876_ _03551_ _03568_ _03574_ _00785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09615_ _00069_ io_in[4] u_cpu.rf_ram.memory\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06827_ u_cpu.rf_ram.memory\[63\]\[5\] _02972_ _02978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06542__A2 _02812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10245__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09546_ u_cpu.rf_ram.memory\[23\]\[1\] _04674_ _04676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08819__A1 _03812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06758_ _02742_ _02934_ _02936_ _00304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05709_ _02188_ _02190_ _02192_ _02194_ _01426_ _02195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__08295__A2 _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09477_ _04637_ _01323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06689_ _02587_ u_cpu.rf_ram.memory\[6\]\[3\] _02894_ _02898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_54_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08428_ _03991_ _03992_ _03997_ _00914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10395__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08359_ u_arbiter.i_wb_cpu_rdt\[24\] u_arbiter.i_wb_cpu_rdt\[8\] _01437_ _03935_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_109_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06058__A1 _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05805__A1 _01553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10321_ _00754_ io_in[4] u_cpu.rf_ram.memory\[34\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09547__A2 _04674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10252_ _00685_ io_in[4] u_cpu.rf_ram.memory\[38\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07558__A1 _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05820__A4 u_cpu.cpu.state.o_cnt_r\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10183_ _00629_ io_in[4] u_cpu.rf_ram.memory\[22\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06230__A1 _01386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05664__S0 _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06781__A2 _02944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07730__A1 _01428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06533__A2 _02801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10738__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08286__A2 _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06297__A1 _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09235__A1 _02577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10888__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05111__I _01547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10519_ _00952_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09538__A2 _04664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10118__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08210__A2 _03800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06221__A1 _02497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05024__A2 _01457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05655__S0 _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05991_ u_cpu.cpu.immdec.imm11_7\[1\] u_cpu.cpu.immdec.imm11_7\[2\] u_cpu.cpu.immdec.imm11_7\[3\]
+ u_cpu.cpu.immdec.imm11_7\[0\] _02452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_38_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10268__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07730_ _01428_ _03451_ _03484_ _03485_ _00727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_04942_ u_cpu.cpu.ctrl.o_ibus_adr\[7\] _01455_ _01459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_37_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05407__S0 _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07661_ u_cpu.rf_ram.memory\[36\]\[3\] _03442_ _03446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_04873_ _01398_ _01399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07721__A1 _03353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06524__A2 _02801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09400_ _04594_ _04595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_77_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06612_ _02738_ _02854_ _02855_ _00239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_19_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07592_ _03353_ _03402_ _03407_ _00667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_18_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09331_ _04474_ _04546_ _04549_ _01265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06543_ u_cpu.rf_ram.memory\[40\]\[3\] _02812_ _02816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06288__A1 _02512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09262_ u_cpu.rf_ram.memory\[85\]\[4\] _04506_ _04511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06474_ _02311_ _02448_ _02367_ _02770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08213_ _03774_ _03781_ _03811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05425_ _01601_ _01913_ _01626_ _01914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_18_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09193_ _04469_ _04470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08029__A2 _02781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09226__A1 _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05356_ _01553_ _01845_ _01654_ _01846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08144_ u_arbiter.i_wb_cpu_rdt\[7\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[7\]
+ _01434_ _03744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07788__A1 _03347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08075_ u_arbiter.i_wb_cpu_rdt\[15\] _03669_ _03678_ u_arbiter.i_wb_cpu_dbus_dat\[15\]
+ _03700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05287_ u_cpu.rf_ram.memory\[132\]\[1\] u_cpu.rf_ram.memory\[133\]\[1\] u_cpu.rf_ram.memory\[134\]\[1\]
+ u_cpu.rf_ram.memory\[135\]\[1\] _01687_ _01688_ _01778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07149__S _03148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09529__A2 _04664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07026_ u_cpu.rf_ram.memory\[53\]\[6\] _03081_ _03088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08201__A2 u_arbiter.i_wb_cpu_rdt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06212__A1 _02475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07260__I0 _02590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05646__S0 _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08977_ u_cpu.rf_ram.memory\[101\]\[0\] _04349_ _04350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07960__A1 _03547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06763__A2 _02934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09903__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07928_ _03551_ _03596_ _03602_ _00809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07859_ u_cpu.rf_ram.memory\[118\]\[6\] _03558_ _03565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06515__A2 _02791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10870_ _01299_ io_in[4] u_cpu.rf_ram.memory\[26\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09529_ _04472_ _04664_ _04666_ _01346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05640__B _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09217__A1 _02684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07059__S _03100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05254__A2 _01744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10304_ _00737_ io_in[4] u_cpu.rf_ram.memory\[92\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06451__A1 _02561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10235_ _00675_ io_in[4] u_cpu.rf_ram.memory\[123\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10410__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05637__S0 _01687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10166_ _00612_ io_in[4] u_cpu.rf_ram.memory\[130\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09583__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07951__A1 _02682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10097_ _00543_ io_in[4] u_cpu.rf_ram.memory\[137\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10560__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07703__A1 _03353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06506__A2 _02791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08751__I0 _02581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05106__I _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08259__A2 _03800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09456__A1 _04468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10999_ _10999_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_90_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05580__I3 u_cpu.rf_ram.memory\[59\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05210_ u_cpu.rf_ram.memory\[0\]\[1\] u_cpu.rf_ram.memory\[1\]\[1\] u_cpu.rf_ram.memory\[2\]\[1\]
+ u_cpu.rf_ram.memory\[3\]\[1\] _01556_ _01557_ _01701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_06190_ _02599_ u_cpu.rf_ram.memory\[1\]\[7\] _02578_ _02600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__05493__A2 _01980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05141_ _01597_ _01632_ _01633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08431__A2 _03809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05072_ _01407_ _01414_ _01564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05709__C _01426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08900_ _04296_ _04299_ _04307_ _01076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06993__A2 _03061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09926__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09880_ _00334_ io_in[4] u_cpu.rf_ram.memory\[63\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10090__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05628__S0 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08831_ _04261_ _04263_ _03797_ _04264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07942__A1 _03547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10903__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06745__A2 _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08762_ _04215_ _01030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05974_ _02309_ u_cpu.cpu.bufreg.c_r _02437_ _02438_ _02439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_66_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07713_ _03343_ _03475_ _03476_ _00719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04925_ u_cpu.cpu.ctrl.o_ibus_adr\[3\] _01439_ _01446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_66_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08693_ _04176_ _01000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_93_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07644_ _03351_ _03432_ _03436_ _00690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04856_ u_cpu.cpu.decode.op21 _01380_ _01381_ _01382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05800__S0 _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07575_ u_cpu.rf_ram.memory\[125\]\[5\] _03392_ _03398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09314_ u_cpu.rf_ram.memory\[111\]\[3\] _04536_ _04540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04855__I u_cpu.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05460__B _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06526_ u_cpu.rf_ram.memory\[17\]\[4\] _02801_ _02806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[61\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09245_ _04501_ _01227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06457_ _02759_ _00180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08670__A2 _04155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05323__I3 u_cpu.rf_ram.memory\[39\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05408_ _01609_ _01896_ _01897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05484__A2 _01971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09176_ _04280_ _04459_ _04460_ _01199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06388_ _02612_ _02684_ _02717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08127_ _03543_ _03731_ _03733_ _00877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05339_ u_cpu.rf_ram.memory\[124\]\[2\] u_cpu.rf_ram.memory\[125\]\[2\] u_cpu.rf_ram.memory\[126\]\[2\]
+ u_cpu.rf_ram.memory\[127\]\[2\] _01545_ _01642_ _01829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_107_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10433__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07481__I0 _02599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08058_ u_arbiter.i_wb_cpu_rdt\[9\] _03669_ _03678_ u_arbiter.i_wb_cpu_dbus_dat\[9\]
+ _03689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_135_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06984__A2 _03061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07009_ _02967_ _03071_ _03078_ _00413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08186__A1 _03776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05619__S0 _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10020_ _00466_ io_in[4] u_cpu.rf_ram.memory\[140\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10583__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07933__A1 _02638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08011__B _02781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08489__A2 _03776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10922_ _01351_ io_in[4] u_cpu.rf_ram.memory\[89\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10853_ _01282_ io_in[4] u_cpu.cpu.genblk3.csr.mcause3_0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09438__A1 _04468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10784_ _01213_ io_in[4] u_cpu.rf_ram.memory\[84\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06672__A1 _02746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09949__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[48\] u_scanchain_local.module_data_in\[47\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[10\] u_scanchain_local.clk u_scanchain_local.module_data_in\[48\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_114_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06424__A1 _02517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05227__A2 _01717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10926__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06975__A2 _03051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08177__A1 _01435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10218_ _00664_ io_in[4] u_cpu.rf_ram.memory\[124\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07924__A1 _03547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06727__A2 _02914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10149_ _00595_ io_in[4] u_cpu.rf_ram.memory\[132\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08724__I0 _02381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05690_ _02169_ _02171_ _02173_ _02175_ _01628_ _02176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_62_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07252__S _03215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10306__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05163__A1 _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05280__B _01402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07360_ u_cpu.rf_ram.memory\[135\]\[0\] _03275_ _03276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04910__A1 u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06311_ _02639_ _02671_ _02672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07291_ _03161_ _03235_ _03237_ _00536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08652__A2 _04145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10456__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09030_ _04378_ _04379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06242_ u_cpu.rf_ram.memory\[78\]\[3\] _02628_ _02632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05466__A2 _01954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06663__A1 _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06173_ _02586_ _02587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08404__A2 _03796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05218__A2 _01708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05124_ _01547_ _01616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05769__A3 _02234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06966__A2 _03051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05055_ u_cpu.raddr\[1\] _01547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09932_ _00386_ io_in[4] u_cpu.rf_ram.memory\[57\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__04977__A1 u_cpu.cpu.ctrl.o_ibus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09863_ _00317_ io_in[4] u_cpu.rf_ram.memory\[64\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07915__A1 _02612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08963__I0 u_arbiter.i_wb_cpu_rdt\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08814_ _03762_ _03778_ _04248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09794_ _00248_ io_in[4] u_cpu.rf_ram.memory\[74\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07391__A2 _03285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08745_ _03553_ _04199_ _04206_ _01022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05174__C _01426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05957_ _01403_ _02416_ _02427_ _00011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_54_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04908_ u_arbiter.i_wb_cpu_ibus_adr\[0\] _01431_ _01432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_27_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08676_ u_cpu.cpu.ctrl.o_ibus_adr\[9\] _04155_ _04157_ u_cpu.cpu.ctrl.o_ibus_adr\[10\]
+ _04167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_53_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05888_ u_cpu.cpu.state.init_done _02367_ _02369_ _02370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_53_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08340__A1 _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07627_ u_cpu.rf_ram.memory\[38\]\[4\] _03422_ _03427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04839_ u_cpu.rf_ram_if.rcnt\[2\] u_cpu.rf_ram_if.rcnt\[1\] _01366_ _01367_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_42_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08891__A2 _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07558_ _03355_ _03382_ _03388_ _00652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__04901__A1 _01406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06509_ _02748_ _02791_ _02796_ _00195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07489_ u_cpu.rf_ram.memory\[22\]\[1\] _03345_ _03348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08643__A2 _04145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06654__A1 _02746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09228_ _04478_ _04487_ _04492_ _01219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_6_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10949__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09159_ u_cpu.rf_ram.memory\[108\]\[1\] _04449_ _04451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05209__A2 _01699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06957__A2 _03041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04968__A1 _01445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08159__A1 _02765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11052_ _11052_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_89_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06709__A2 _02904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10003_ _00449_ io_in[4] u_cpu.rf_ram.memory\[142\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05068__S1 _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05365__B _01417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07382__A2 _03285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10329__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08168__S _01436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09621__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07072__S _03109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07134__A2 _03139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10905_ _01334_ io_in[4] u_cpu.rf_ram.memory\[98\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08882__A2 _04282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10479__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05696__A2 _02181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10836_ _01265_ io_in[4] u_cpu.rf_ram.memory\[87\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10767_ _01196_ io_in[4] u_cpu.rf_ram.memory\[108\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09771__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06645__A1 _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10698_ _01127_ io_in[4] u_cpu.rf_ram.memory\[103\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08398__A1 _03743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08398__B2 _03831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05259__C _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06948__A2 _03041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05620__A2 _02106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08945__I0 u_arbiter.i_wb_cpu_rdt\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05059__S1 _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06860_ _02961_ _02992_ _02996_ _00346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07373__A2 _03275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05811_ u_cpu.rf_ram.memory\[140\]\[7\] u_cpu.rf_ram.memory\[141\]\[7\] u_cpu.rf_ram.memory\[142\]\[7\]
+ u_cpu.rf_ram.memory\[143\]\[7\] _01680_ _01681_ _02296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_83_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06791_ _02954_ _02955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08530_ u_cpu.rf_ram.memory\[32\]\[1\] _04084_ _04086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05742_ _01570_ _02226_ _02227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07125__A2 _03139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08461_ _03778_ _03786_ _04025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05673_ u_cpu.rf_ram.memory\[44\]\[6\] u_cpu.rf_ram.memory\[45\]\[6\] u_cpu.rf_ram.memory\[46\]\[6\]
+ u_cpu.rf_ram.memory\[47\]\[6\] _01615_ _01616_ _02159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08873__A2 _04282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07676__A3 _03454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07412_ _02561_ _02832_ _03304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05231__S1 _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06884__A1 _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08392_ _03812_ _03961_ _03962_ _03964_ _03965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_32_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08086__B1 _03678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07343_ _03157_ _03265_ _03266_ _00559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08625__A2 _02394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06636__A1 _02746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07274_ u_cpu.rf_ram.memory\[138\]\[2\] _03225_ _03228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09013_ u_cpu.rf_ram.memory\[103\]\[0\] _04369_ _04370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06225_ _02507_ _02614_ _02620_ _00087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08389__A1 _03761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08389__B2 _03788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06156_ _02572_ _02573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09050__A2 _04389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06939__A2 _03031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05107_ u_cpu.rf_ram.memory\[60\]\[0\] u_cpu.rf_ram.memory\[61\]\[0\] u_cpu.rf_ram.memory\[62\]\[0\]
+ u_cpu.rf_ram.memory\[63\]\[0\] _01598_ _01573_ _01599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_132_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05298__S1 _01557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06087_ _02492_ _02530_ _02533_ _00036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05964__I u_cpu.cpu.bufreg.lsb\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09915_ _00369_ io_in[4] u_cpu.rf_ram.memory\[5\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05038_ u_cpu.cpu.ctrl.o_ibus_adr\[29\] u_cpu.cpu.ctrl.o_ibus_adr\[28\] u_cpu.cpu.ctrl.o_ibus_adr\[27\]
+ _01523_ _01532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_58_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09846_ _00300_ io_in[4] u_cpu.rf_ram.memory\[66\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09644__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07364__A2 _03275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08561__A1 _03555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09777_ _00231_ io_in[4] u_cpu.rf_ram.memory\[139\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06989_ _02965_ _03061_ _03067_ _00404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08728_ _04196_ _01015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05470__S1 _01557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10621__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07116__A2 _03129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08659_ _04158_ _00984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_14_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09794__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08864__A2 _04282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05222__S1 _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10621_ _01050_ io_in[4] u_cpu.cpu.immdec.imm11_7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10771__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06627__A1 _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10552_ _00024_ io_in[4] u_cpu.cpu.ctrl.pc_plus_offset_cy_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10483_ _00916_ io_in[4] u_cpu.cpu.immdec.imm19_12_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10001__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09041__A2 _04379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11104_ _11104_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_111_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10151__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11035_ _11035_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__05095__B _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07355__A2 _03265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05461__S1 _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08304__A1 _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07107__A2 _03129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05542__C _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06166__I0 _02581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08855__A2 _04271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05669__A2 _02154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05213__S1 _01574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06866__A1 _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10819_ _01248_ io_in[4] u_cpu.rf_ram.memory\[86\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06618__A1 _02746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09280__A2 _04516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07291__A1 _03161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06094__A2 _02530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06010_ _02466_ _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09032__A2 _04379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07043__A1 _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07594__A2 _03402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09667__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08791__A1 _03547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07961_ u_cpu.rf_ram.memory\[115\]\[4\] _03616_ _03621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[34\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09700_ _00154_ io_in[4] u_cpu.rf_ram.memory\[48\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06912_ _02587_ u_cpu.rf_ram.memory\[5\]\[3\] _03021_ _03025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07892_ _02593_ u_cpu.rf_ram.memory\[8\]\[5\] _03577_ _03583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10644__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08543__A1 _03555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07346__A2 _03265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09631_ _00085_ io_in[4] u_cpu.rf_ram.memory\[80\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06843_ u_cpu.rf_ram.memory\[62\]\[4\] _02982_ _02987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05452__S1 _01549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09562_ _04155_ _04683_ _04684_ _01361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06774_ _02738_ _02944_ _02945_ _00311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09099__A2 _04409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[49\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08513_ _01375_ u_cpu.cpu.immdec.imm24_20\[0\] _04073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05725_ u_cpu.rf_ram.memory\[128\]\[6\] u_cpu.rf_ram.memory\[129\]\[6\] u_cpu.rf_ram.memory\[130\]\[6\]
+ u_cpu.rf_ram.memory\[131\]\[6\] _01572_ _01688_ _02211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_70_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09493_ _04472_ _04644_ _04646_ _01330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10794__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08846__A2 _04271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08444_ _04010_ _04011_ _04012_ _03798_ _00915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__05204__S1 _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05904__I0 u_arbiter.i_wb_cpu_dbus_dat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05656_ _01562_ _02141_ _01582_ _02142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08375_ _02765_ u_arbiter.i_wb_cpu_rdt\[25\] _03950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05587_ u_cpu.rf_ram.memory\[36\]\[5\] u_cpu.rf_ram.memory\[37\]\[5\] u_cpu.rf_ram.memory\[38\]\[5\]
+ u_cpu.rf_ram.memory\[39\]\[5\] _01619_ _01620_ _02074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_23_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10024__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06609__A1 _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07326_ u_cpu.rf_ram.memory\[49\]\[1\] _03255_ _03257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06085__A2 _02530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07257_ _03218_ _00521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06208_ _02610_ _00080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09023__A2 _04369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07188_ _03165_ _03176_ _03180_ _00490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10174__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06139_ u_cpu.rf_ram.memory\[20\]\[0\] _02563_ _02564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07585__A2 _03402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08782__A1 _02475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05140__S0 _01619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05691__S1 _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07337__A2 _03255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05348__A1 _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09829_ _00283_ io_in[4] u_cpu.rf_ram.memory\[68\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05643__B _02129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05443__S1 _01652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08837__A2 _03798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06848__A1 _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07896__I0 _02599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05520__A1 _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10604_ _01033_ io_in[4] u_cpu.rf_ram.memory\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09262__A2 _04506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10517__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10535_ _00968_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07273__A1 _03161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10466_ _00899_ io_in[4] u_cpu.rf_ram.memory\[114\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09014__A2 _04369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[30\] u_arbiter.i_wb_cpu_rdt\[27\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[24\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__07025__A1 _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09565__A3 u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10397_ _00830_ io_in[4] u_cpu.rf_ram.memory\[116\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10667__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07576__A2 _03392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05682__S1 _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05109__I _01540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07328__A2 _03255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11018_ _11018_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_38_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06000__A2 _01386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05045__S _01431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10047__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05510_ u_cpu.rf_ram.memory\[100\]\[4\] u_cpu.rf_ram.memory\[101\]\[4\] u_cpu.rf_ram.memory\[102\]\[4\]
+ u_cpu.rf_ram.memory\[103\]\[4\] _01577_ _01549_ _01998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_06490_ u_cpu.rf_ram_if.rcnt\[2\] u_cpu.rf_ram_if.rcnt\[1\] u_cpu.rf_ram_if.rcnt\[0\]
+ _02785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_2690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07260__S _03215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05441_ u_cpu.rf_ram.memory\[80\]\[3\] u_cpu.rf_ram.memory\[81\]\[3\] u_cpu.rf_ram.memory\[82\]\[3\]
+ u_cpu.rf_ram.memory\[83\]\[3\] _01590_ _01642_ _01930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_21_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05511__A1 _01636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08160_ _01435_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[3\] _03760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05372_ _01684_ _01861_ _01582_ _01862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10197__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07111_ _02963_ _03129_ _03134_ _00459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08091_ u_arbiter.i_wb_cpu_rdt\[21\] _03653_ _03654_ u_arbiter.i_wb_cpu_dbus_dat\[21\]
+ _03676_ u_arbiter.i_wb_cpu_dbus_dat\[22\] _03710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_109_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07042_ u_cpu.rf_ram.memory\[52\]\[5\] _03091_ _03097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09005__A2 _04359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05728__B _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07567__A2 _03392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[18\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08993_ _02893_ _04197_ _04358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07944_ _03549_ _03606_ _03611_ _00816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05673__S1 _01616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07319__A2 _03245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07875_ u_cpu.rf_ram.memory\[121\]\[5\] _03568_ _03574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09614_ _00068_ io_in[4] u_cpu.rf_ram.memory\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06826_ _02963_ _02972_ _02977_ _00331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__04858__I u_cpu.cpu.genblk3.csr.o_new_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09545_ _04468_ _04674_ _04675_ _01353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06757_ u_cpu.rf_ram.memory\[65\]\[1\] _02934_ _02936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05708_ _01614_ _02193_ _01654_ _02194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_19_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09476_ _02584_ u_cpu.rf_ram.memory\[0\]\[2\] _04634_ _04637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06688_ _02897_ _00273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_58_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09492__A2 _04644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08493__C _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08427_ u_cpu.cpu.immdec.imm7 _02438_ _03956_ _03996_ _03997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_24_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05502__A1 _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05639_ u_cpu.rf_ram.memory\[132\]\[5\] u_cpu.rf_ram.memory\[133\]\[5\] u_cpu.rf_ram.memory\[134\]\[5\]
+ u_cpu.rf_ram.memory\[135\]\[5\] _01687_ _01688_ _02126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08358_ _03741_ _03786_ _03820_ _03756_ _03859_ _03934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__09832__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06058__A2 u_cpu.rf_ram_if.wdata1_r\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07309_ _03161_ _03245_ _03247_ _00544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08289_ _02469_ _02821_ _03878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10320_ _00753_ io_in[4] u_cpu.rf_ram.memory\[34\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07007__A1 _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10251_ _00684_ io_in[4] u_cpu.rf_ram.memory\[38\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09982__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07558__A2 _03382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05357__C _01426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10182_ _00628_ io_in[4] u_cpu.rf_ram.memory\[22\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05664__S1 _01548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08507__A1 _03741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09180__A1 _04286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07080__S _03109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06297__A2 _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[32\]_D u_arbiter.i_wb_cpu_rdt\[29\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09235__A2 _02638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07246__A1 _03169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07797__A2 _03520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10518_ _00951_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10449_ _00882_ io_in[4] u_cpu.rf_ram.memory\[113\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05548__B _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07549__A2 _03382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08210__A3 _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06221__A2 _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05655__S1 _01580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05990_ _01387_ _02433_ u_cpu.cpu.o_wen1 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04941_ _01454_ _01456_ _01458_ u_arbiter.o_wb_cpu_adr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09705__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05407__S1 _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07660_ _03349_ _03442_ _03445_ _00697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04872_ _01397_ _01398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_92_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07721__A2 _03475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06611_ u_cpu.rf_ram.memory\[77\]\[0\] _02854_ _02855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07591_ u_cpu.rf_ram.memory\[124\]\[4\] _03402_ _03407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09330_ u_cpu.rf_ram.memory\[87\]\[2\] _04546_ _04549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06542_ _02744_ _02812_ _02815_ _00209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09855__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06288__A2 _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09261_ _04476_ _04506_ _04510_ _01234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06473_ _01428_ _02769_ _00186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08682__B1 _04157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08212_ _03803_ _03809_ _03810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05424_ u_cpu.rf_ram.memory\[96\]\[3\] u_cpu.rf_ram.memory\[97\]\[3\] u_cpu.rf_ram.memory\[98\]\[3\]
+ u_cpu.rf_ram.memory\[99\]\[3\] _01602_ _01579_ _01913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10832__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09192_ _02475_ _02561_ _04469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_u_scanchain_local.scan_flop\[23\]_D u_arbiter.i_wb_cpu_rdt\[20\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09226__A2 _04487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08143_ u_arbiter.i_wb_cpu_rdt\[9\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[9\]
+ _01435_ _03743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05355_ u_cpu.rf_ram.memory\[84\]\[2\] u_cpu.rf_ram.memory\[85\]\[2\] u_cpu.rf_ram.memory\[86\]\[2\]
+ u_cpu.rf_ram.memory\[87\]\[2\] _01555_ _01652_ _01845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07788__A2 _03520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08074_ u_arbiter.i_wb_cpu_dbus_dat\[16\] _03683_ _03699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05343__S0 _01619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05286_ _01399_ _01776_ _01777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05799__A1 _01667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07025_ _02965_ _03081_ _03087_ _00420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08737__A1 _03545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06212__A2 _02612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10212__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05646__S1 _01557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08976_ _04348_ _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07960__A2 _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07927_ u_cpu.rf_ram.memory\[112\]\[5\] _03596_ _03602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05971__A1 _02436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09162__A1 _04286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07858_ _03551_ _03558_ _03564_ _00777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07712__A2 _03475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10362__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06809_ _02511_ _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07789_ u_cpu.rf_ram.memory\[34\]\[2\] _03520_ _03523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09528_ u_cpu.rf_ram.memory\[89\]\[1\] _04664_ _04666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09465__A2 _04625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06279__A2 _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09459_ u_cpu.rf_ram.memory\[24\]\[2\] _04625_ _04628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[14\]_D u_arbiter.i_wb_cpu_rdt\[11\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09217__A2 _02706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07228__A1 _03169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07779__A2 _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05334__S0 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10303_ _00736_ io_in[4] u_cpu.rf_ram.memory\[92\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06451__A2 _02577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05368__B _01402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10234_ _00674_ io_in[4] u_cpu.rf_ram.memory\[123\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06043__I _02496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09728__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05637__S1 _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10165_ _00611_ io_in[4] u_cpu.rf_ram.memory\[130\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07951__A2 _02821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10096_ _00542_ io_in[4] u_cpu.rf_ram.memory\[39\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10705__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09878__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07703__A2 _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08900__A1 _04296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10855__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10998_ _10998_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__09456__A2 _04625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08664__B1 _04157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05122__I _01397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05140_ u_cpu.rf_ram.memory\[108\]\[0\] u_cpu.rf_ram.memory\[109\]\[0\] u_cpu.rf_ram.memory\[110\]\[0\]
+ u_cpu.rf_ram.memory\[111\]\[0\] _01619_ _01620_ _01632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_144_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05325__S0 _01623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05071_ u_cpu.rf_ram.memory\[0\]\[0\] u_cpu.rf_ram.memory\[1\]\[0\] u_cpu.rf_ram.memory\[2\]\[0\]
+ u_cpu.rf_ram.memory\[3\]\[0\] _01556_ _01557_ _01563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10235__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08195__A2 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09392__A1 _04191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05628__S1 _01549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08830_ _02525_ _04236_ _04262_ _04263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_44_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07942__A2 _03606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10385__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08761_ _02596_ u_cpu.rf_ram.memory\[3\]\[6\] _04208_ _04215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05973_ _01374_ _02383_ _02438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05953__A1 _01403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09144__A1 _04286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07712_ u_cpu.rf_ram.memory\[90\]\[0\] _03475_ _03476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_04924_ _01442_ _01445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08692_ u_cpu.cpu.ctrl.o_ibus_adr\[16\] _04173_ _04175_ u_cpu.cpu.ctrl.o_ibus_adr\[17\]
+ _04176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_26_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07643_ u_cpu.rf_ram.memory\[37\]\[3\] _03432_ _03436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04855_ u_cpu.cpu.decode.co_ebreak _01381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07574_ _03353_ _03392_ _03397_ _00659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05800__S1 _01652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09447__A2 _04615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09313_ _04474_ _04536_ _04539_ _01257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06525_ _02746_ _02801_ _02805_ _00202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09244_ _02590_ u_cpu.rf_ram.memory\[10\]\[4\] _04496_ _04501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06456_ _02584_ u_cpu.rf_ram.memory\[4\]\[2\] _02756_ _02759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06130__A1 _02507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05407_ u_cpu.rf_ram.memory\[40\]\[3\] u_cpu.rf_ram.memory\[41\]\[3\] u_cpu.rf_ram.memory\[42\]\[3\]
+ u_cpu.rf_ram.memory\[43\]\[3\] _01545_ _01611_ _01896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09175_ u_cpu.rf_ram.memory\[69\]\[0\] _04459_ _04460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06387_ _02517_ _02708_ _02716_ _00153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08126_ u_cpu.rf_ram.memory\[113\]\[1\] _03731_ _03733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05338_ _01821_ _01823_ _01825_ _01827_ _01628_ _01828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_108_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05316__S0 _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07630__A1 _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08057_ u_arbiter.i_wb_cpu_dbus_dat\[10\] _03683_ _03688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05269_ _01753_ _01755_ _01757_ _01759_ _01426_ _01760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_116_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07008_ u_cpu.rf_ram.memory\[54\]\[6\] _03071_ _03078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04995__A2 _01442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10728__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08186__A2 _03785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08499__B _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05619__S1 _01652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07933__A2 _02821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08959_ u_arbiter.i_wb_cpu_rdt\[24\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[8\]
+ _04331_ _04340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__05944__A1 _02321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10878__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10921_ _01350_ io_in[4] u_cpu.rf_ram.memory\[89\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07697__A1 _03347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05651__B _01565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10852_ _01281_ io_in[4] u_cpu.cpu.genblk3.csr.mcause3_0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09438__A2 _04615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10108__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10783_ _01212_ io_in[4] u_cpu.rf_ram.memory\[84\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06672__A2 _02884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10258__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05307__S0 _01578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06424__A2 _02729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10217_ _00663_ io_in[4] u_cpu.rf_ram.memory\[124\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07924__A2 _03596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10148_ _00594_ io_in[4] u_cpu.rf_ram.memory\[132\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05935__A1 _02321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09126__A1 _04286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10079_ _00525_ io_in[4] u_cpu.rf_ram.memory\[14\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05117__I _01540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08724__I1 _02406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06360__A1 _02497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09429__A2 _04605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08488__I0 u_arbiter.i_wb_cpu_rdt\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04910__A2 _01431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06310_ _02560_ _02624_ _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07290_ u_cpu.rf_ram.memory\[39\]\[1\] _03235_ _03237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06112__A1 _02507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06241_ _02492_ _02628_ _02631_ _00092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07860__A1 _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06663__A2 _02706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06172_ u_cpu.rf_ram_if.wdata0_r\[3\] u_cpu.rf_ram_if.wdata1_r\[3\] _02478_ _02586_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_102_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08404__A3 _03947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05123_ _01543_ _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07612__A1 _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06415__A2 _02729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05054_ _01545_ _01546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09931_ _00385_ io_in[4] u_cpu.rf_ram.memory\[57\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09365__A1 _01385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09862_ _00316_ io_in[4] u_cpu.rf_ram.memory\[64\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07915__A2 _02821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08813_ _04245_ _04247_ _01049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05926__A1 _01374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09793_ _00247_ io_in[4] u_cpu.rf_ram.memory\[74\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08744_ u_cpu.rf_ram.memory\[109\]\[6\] _04199_ _04206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05956_ u_cpu.rf_ram_if.rdata0\[4\] _01403_ _02427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_04907_ _01430_ _01431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08675_ _04166_ _00992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__07679__A1 u_cpu.cpu.mem_bytecnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05887_ u_cpu.cpu.state.stage_two_req _02368_ _02369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05471__B _01417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08340__A2 _03914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07626_ _03351_ _03422_ _03426_ _00682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04838_ u_cpu.rf_ram_if.rcnt\[0\] _01366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06351__A1 _02639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05785__S0 _01623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07557_ u_cpu.rf_ram.memory\[126\]\[5\] _03382_ _03388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__04901__A2 _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10400__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06508_ u_cpu.rf_ram.memory\[16\]\[4\] _02791_ _02796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07488_ _02486_ _03347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07151__I0 _02599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09573__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06654__A2 _02874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09227_ u_cpu.rf_ram.memory\[59\]\[4\] _04487_ _04492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06439_ _02501_ _02748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09158_ _04280_ _04449_ _04450_ _01191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08109_ u_arbiter.i_wb_cpu_rdt\[27\] _03653_ _03654_ u_arbiter.i_wb_cpu_dbus_dat\[27\]
+ _03722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10550__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09089_ u_cpu.rf_ram.memory\[105\]\[2\] _04409_ _04412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08159__A2 u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11051_ _11051_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_107_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10002_ _00448_ io_in[4] u_cpu.rf_ram.memory\[142\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05917__A1 _02394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09108__A1 _04286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06590__A1 _02754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10904_ _01333_ io_in[4] u_cpu.rf_ram.memory\[98\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05776__S0 _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10835_ _01264_ io_in[4] u_cpu.rf_ram.memory\[87\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06893__A2 _03012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09916__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10080__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10766_ _01195_ io_in[4] u_cpu.rf_ram.memory\[108\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[60\] u_scanchain_local.module_data_in\[59\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[22\] u_scanchain_local.clk u_scanchain_local.module_data_in\[60\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_40_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06645__A2 _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10697_ _01126_ io_in[4] u_cpu.rf_ram.memory\[102\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08398__A2 _03786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09347__A1 _04472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[51\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05908__A1 _01373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05810_ _01399_ _02294_ _02295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06790_ _02528_ _02660_ _02954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08359__S _01437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05741_ u_cpu.rf_ram.memory\[20\]\[7\] u_cpu.rf_ram.memory\[21\]\[7\] u_cpu.rf_ram.memory\[22\]\[7\]
+ u_cpu.rf_ram.memory\[23\]\[7\] _01572_ _01574_ _02226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_82_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10423__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08460_ _03973_ _03988_ _03801_ _04024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05672_ _01609_ _02157_ _02158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06184__I1 u_cpu.rf_ram_if.wdata1_r\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07411_ _03173_ _03295_ _03303_ _00590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_17_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08391_ _03788_ _03896_ _03963_ _03779_ _03851_ _03964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_51_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09596__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06884__A2 _03002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04895__A1 _01419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07342_ u_cpu.rf_ram.memory\[136\]\[0\] _03265_ _03266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05519__S0 _01619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10573__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07273_ _03161_ _03225_ _03227_ _00528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06636__A2 _02864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09012_ _04368_ _04369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06224_ u_cpu.rf_ram.memory\[80\]\[5\] _02614_ _02620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08389__A2 _03860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06155_ u_cpu.rf_ram_if.wdata0_r\[0\] u_cpu.rf_ram_if.wdata1_r\[0\] _02478_ _02572_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05106_ _01544_ _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06086_ u_cpu.rf_ram.memory\[21\]\[2\] _02530_ _02533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09914_ _00368_ io_in[4] u_cpu.rf_ram.memory\[5\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05037_ _01443_ _01530_ _01531_ u_arbiter.o_wb_cpu_adr\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_63_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08010__A1 _03648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09845_ _00299_ io_in[4] u_cpu.rf_ram.memory\[66\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05185__C _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08561__A2 _04094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09776_ _00230_ io_in[4] u_cpu.rf_ram.memory\[129\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_101_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05980__I _02372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06988_ u_cpu.rf_ram.memory\[55\]\[5\] _03061_ _03067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08727_ u_cpu.cpu.ctrl.o_ibus_adr\[31\] _04154_ _04175_ _04195_ _04196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05939_ _02320_ u_cpu.rf_ram_if.rdata1\[3\] _02417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_2_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09939__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06324__A1 _02507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08658_ u_arbiter.i_wb_cpu_ibus_adr\[0\] _04155_ _04157_ u_arbiter.i_wb_cpu_ibus_adr\[1\]
+ _04158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_15_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07901__S _03586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07609_ u_cpu.rf_ram.memory\[123\]\[4\] _03412_ _03417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10916__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06875__A2 _03002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08589_ u_arbiter.i_wb_cpu_dbus_adr\[15\] u_arbiter.i_wb_cpu_dbus_adr\[14\] _04115_
+ _04117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10620_ _01049_ io_in[4] u_cpu.cpu.immdec.imm11_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10551_ _00983_ io_in[4] u_cpu.rf_ram.memory\[30\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06627__A2 _02638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10482_ _00915_ io_in[4] u_cpu.cpu.immdec.imm7 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11103_ _11103_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__09329__A1 _04472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05376__B _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11034_ _11034_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_104_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08552__A2 _04094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10446__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06563__A1 _02746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05366__A2 _01851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09501__A1 _04480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08304__A2 _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10596__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06866__A2 _02992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10818_ _01247_ io_in[4] u_cpu.rf_ram.memory\[86\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06618__A2 _02854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10749_ _01178_ io_in[4] u_cpu.rf_ram.memory\[107\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07291__A2 _03235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07258__S _03215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08240__A1 _02333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06162__S _02578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07043__A2 _03091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08791__A2 _04227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07960_ _03547_ _03616_ _03620_ _00823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06911_ _03024_ _00369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07891_ _03582_ _00792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08543__A2 _04084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09630_ _00084_ io_in[4] u_cpu.rf_ram.memory\[80\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06842_ _02961_ _02982_ _02986_ _00338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06554__A1 _02602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05357__A2 _01842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09561_ u_cpu.cpu.state.ibus_cyc _04683_ _04684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06773_ u_cpu.rf_ram.memory\[64\]\[0\] _02944_ _02945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10939__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08512_ _03741_ _04027_ _04068_ _03791_ _04071_ _04072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_05724_ _01684_ _02209_ _01582_ _02210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09492_ u_cpu.rf_ram.memory\[98\]\[1\] _04644_ _04646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08443_ u_cpu.cpu.immdec.imm7 _02305_ _04012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06857__A2 _02992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05655_ u_cpu.rf_ram.memory\[16\]\[6\] u_cpu.rf_ram.memory\[17\]\[6\] u_cpu.rf_ram.memory\[18\]\[6\]
+ u_cpu.rf_ram.memory\[19\]\[6\] _01556_ _01580_ _02141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_23_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05904__I1 u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04868__A1 u_cpu.cpu.decode.op21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08374_ _03797_ _03948_ _03949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05586_ _01397_ _02072_ _01605_ _02073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_108_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07325_ _03157_ _03255_ _03256_ _00551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07806__A1 _03347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06609__A2 _02660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05817__B1 _02299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07256_ _02584_ u_cpu.rf_ram.memory\[14\]\[2\] _03215_ _03218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07282__A2 _03225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10319__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05293__A1 _01542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06207_ _02596_ u_cpu.rf_ram.memory\[7\]\[6\] _02603_ _02610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09559__A1 _04484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07187_ u_cpu.rf_ram.memory\[73\]\[3\] _03176_ _03180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09611__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06138_ _02562_ _02563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08231__A1 _03767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07034__A2 _03091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08782__A2 _02660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06069_ _02477_ _02517_ _02518_ _00033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10469__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05140__S1 _01620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06793__A1 _02953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09761__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08534__A2 _04084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09828_ _00282_ io_in[4] u_cpu.rf_ram.memory\[68\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05348__A2 _01828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09759_ _00213_ io_in[4] u_cpu.rf_ram.memory\[40\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08298__A1 _03547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06848__A2 _02982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05520__A2 _02007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10603_ _01032_ io_in[4] u_cpu.rf_ram.memory\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08470__A1 _03999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10534_ _00967_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07273__A2 _03225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05284__A1 _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10465_ _00898_ io_in[4] u_cpu.rf_ram.memory\[114\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07078__S _03109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08222__A1 _03741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07025__A2 _03081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10396_ _00829_ io_in[4] u_cpu.rf_ram.memory\[116\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05036__A1 u_arbiter.i_wb_cpu_dbus_adr\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[23\] u_arbiter.i_wb_cpu_rdt\[20\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[17\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_2_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06784__A1 _02750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11017_ _11017_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_93_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05553__C _01404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08289__A1 _02469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06839__A2 _02982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05440_ _01645_ _01928_ _01648_ _01929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_33_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05371_ u_cpu.rf_ram.memory\[140\]\[2\] u_cpu.rf_ram.memory\[141\]\[2\] u_cpu.rf_ram.memory\[142\]\[2\]
+ u_cpu.rf_ram.memory\[143\]\[2\] _01680_ _01681_ _01861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07110_ u_cpu.rf_ram.memory\[141\]\[4\] _03129_ _03134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09634__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08090_ _03708_ _03709_ _00864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08461__A1 _03778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05275__A1 _01667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07041_ _02963_ _03091_ _03096_ _00427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10611__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08213__A1 _03774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07016__A2 _03081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09784__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08992_ _04296_ _04349_ _04357_ _01118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_141_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07943_ u_cpu.rf_ram.memory\[122\]\[4\] _03606_ _03611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10761__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08516__A2 _04016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05744__B _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07874_ _03549_ _03568_ _03573_ _00784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06527__A1 _02748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09613_ _00067_ io_in[4] u_cpu.rf_ram.memory\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06825_ u_cpu.rf_ram.memory\[63\]\[4\] _02972_ _02977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09544_ u_cpu.rf_ram.memory\[23\]\[0\] _04674_ _04675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06756_ _02738_ _02934_ _02935_ _00303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05707_ u_cpu.rf_ram.memory\[84\]\[6\] u_cpu.rf_ram.memory\[85\]\[6\] u_cpu.rf_ram.memory\[86\]\[6\]
+ u_cpu.rf_ram.memory\[87\]\[6\] _01555_ _01652_ _02193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_93_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06687_ _02584_ u_cpu.rf_ram.memory\[6\]\[2\] _02894_ _02897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09475_ _04636_ _01322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_19_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08426_ _03993_ _03994_ _03995_ _02438_ _03996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05638_ _01399_ _02124_ _02125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05502__A2 _01989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10141__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08357_ _03916_ _03931_ _03932_ _03933_ _00907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_05569_ u_cpu.rf_ram.memory\[28\]\[5\] u_cpu.rf_ram.memory\[29\]\[5\] u_cpu.rf_ram.memory\[30\]\[5\]
+ u_cpu.rf_ram.memory\[31\]\[5\] _01572_ _01574_ _02056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_20_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07308_ u_cpu.rf_ram.memory\[137\]\[1\] _03245_ _03247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08288_ _02337_ _03740_ _03877_ _00894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05266__A1 _01609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07239_ u_cpu.rf_ram.memory\[143\]\[2\] _03206_ _03209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10291__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10250_ _00683_ io_in[4] u_cpu.rf_ram.memory\[38\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08204__A1 _03767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07007__A2 _03071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10181_ _00627_ io_in[4] u_cpu.rf_ram.memory\[22\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06766__A1 _02750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08507__A2 _03988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09180__A2 _04459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09657__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[33\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10634__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07246__A2 _03206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10517_ _00950_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_u_scanchain_local.scan_flop\[48\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10448_ _00881_ io_in[4] u_cpu.rf_ram.memory\[113\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05009__A1 _01443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10784__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08746__A2 _04199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10379_ _00812_ io_in[4] u_cpu.rf_ram.memory\[122\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04940_ u_arbiter.i_wb_cpu_dbus_adr\[6\] _01457_ _01458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10014__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06509__A1 _02748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09171__A2 _04449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04871_ _01396_ _01397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07182__A1 _03157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06610_ _02853_ _02854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07590_ _03351_ _03402_ _03406_ _00666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_19_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10164__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06541_ u_cpu.rf_ram.memory\[40\]\[2\] _02812_ _02815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09260_ u_cpu.rf_ram.memory\[85\]\[3\] _04506_ _04510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06472_ u_cpu.cpu.state.genblk1.misalign_trap_sync_r u_cpu.cpu.state.stage_two_req
+ _02768_ _02769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_34_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05496__A1 _01609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05423_ _01636_ _01911_ _01912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08211_ _03776_ _03768_ _03809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09191_ _02481_ _04468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05354_ _01609_ _01843_ _01844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08142_ u_arbiter.i_wb_cpu_rdt\[10\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[10\]
+ _01434_ _03742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09482__I0 _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08434__A1 _03831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07237__A2 _03206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08985__A2 _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08073_ _03698_ _00858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_135_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05739__B _01565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05285_ u_cpu.rf_ram.memory\[128\]\[1\] u_cpu.rf_ram.memory\[129\]\[1\] u_cpu.rf_ram.memory\[130\]\[1\]
+ u_cpu.rf_ram.memory\[131\]\[1\] _01687_ _01688_ _01776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_88_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05343__S1 _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05799__A2 _02283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07024_ u_cpu.rf_ram.memory\[53\]\[5\] _03081_ _03087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08737__A2 _04199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06748__A1 _02750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08975_ _02524_ _04197_ _04348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07926_ _03549_ _03596_ _03601_ _00808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05971__A2 _01431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09162__A2 _04449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07857_ u_cpu.rf_ram.memory\[118\]\[5\] _03558_ _03564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10507__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08370__B1 _03800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06808_ _02965_ _02955_ _02966_ _00324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08277__S _01436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07788_ _03347_ _03520_ _03522_ _00749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09527_ _04468_ _04664_ _04665_ _01345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06739_ u_cpu.rf_ram.memory\[66\]\[1\] _02924_ _02926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10657__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09458_ _04472_ _04625_ _04627_ _01314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05487__A1 _01589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08409_ _03776_ _03851_ _03980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_8_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09389_ _04584_ _04586_ _04587_ _01285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_40_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07228__A2 _03196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05239__B2 _01729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05334__S1 _01549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06987__A1 _02963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08025__B _02774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10302_ _00735_ io_in[4] u_cpu.rf_ram.memory\[92\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10233_ _00673_ io_in[4] u_cpu.rf_ram.memory\[123\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10037__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10164_ _00610_ io_in[4] u_cpu.rf_ram.memory\[130\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07400__A2 _03295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10095_ _00541_ io_in[4] u_cpu.rf_ram.memory\[39\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05962__A2 _01403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10187__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09153__A2 _04439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08361__B1 _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08900__A2 _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05565__I2 u_cpu.rf_ram.memory\[22\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05270__S0 _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[2\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10997_ _10997_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_76_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05478__A1 _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08416__A1 _03742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07219__A2 _03196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05559__B _01417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05325__S1 _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05070_ _01541_ _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05278__C _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07266__S _03215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05089__S0 _01578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06170__S _02578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08760_ _04214_ _01029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05972_ _01374_ u_cpu.cpu.decode.opcode\[1\] _02437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09822__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07711_ _03474_ _03475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09144__A2 _04439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04923_ _01438_ _01440_ _01444_ u_arbiter.o_wb_cpu_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08691_ _04156_ _04175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07642_ _03349_ _03432_ _03435_ _00689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_04854_ u_cpu.cpu.decode.op26 _01380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_53_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06902__A1 _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05261__S0 _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07573_ u_cpu.rf_ram.memory\[125\]\[4\] _03392_ _03397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08104__B1 _03654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09972__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09312_ u_cpu.rf_ram.memory\[111\]\[2\] _04536_ _04539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06524_ u_cpu.rf_ram.memory\[17\]\[3\] _02801_ _02805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07458__A2 _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05469__A1 _01542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09243_ _04500_ _01226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06455_ _02758_ _00179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06130__A2 _02551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08407__A1 _01437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05406_ _01888_ _01890_ _01892_ _01894_ _01607_ _01895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_06386_ u_cpu.rf_ram.memory\[43\]\[7\] _02708_ _02716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09174_ _04458_ _04459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08125_ _03539_ _03731_ _03732_ _00876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05337_ _01601_ _01826_ _01626_ _01827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09080__A1 _04294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05316__S1 _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06969__A1 _02963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05268_ _01553_ _01758_ _01654_ _01759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08056_ _03686_ _03687_ _00852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07630__A2 _03422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07007_ _02965_ _03071_ _03077_ _00412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05199_ u_cpu.rf_ram.memory\[132\]\[0\] u_cpu.rf_ram.memory\[133\]\[0\] u_cpu.rf_ram.memory\[134\]\[0\]
+ u_cpu.rf_ram.memory\[135\]\[0\] _01687_ _01688_ _01691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_143_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07394__A1 _02524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08958_ _04339_ _01102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09135__A2 _04429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07909_ _02593_ u_cpu.rf_ram.memory\[11\]\[5\] _03586_ _03592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08889_ u_cpu.rf_ram.memory\[95\]\[2\] _04299_ _04302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10920_ _01349_ io_in[4] u_cpu.rf_ram.memory\[89\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07697__A2 _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08894__A1 _04290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10851_ _01280_ io_in[4] u_cpu.cpu.genblk3.csr.mcause3_0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10782_ _01211_ io_in[4] u_cpu.rf_ram.memory\[84\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06121__A2 _02551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05307__S1 _01580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07621__A2 _03422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05632__A1 _02099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09845__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10216_ _00662_ io_in[4] u_cpu.rf_ram.memory\[125\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09374__A2 _04568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07385__A1 _03165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10147_ _00593_ io_in[4] u_cpu.rf_ram.memory\[132\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10822__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09126__A2 _04429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10078_ _00524_ io_in[4] u_cpu.rf_ram.memory\[14\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09995__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05699__A1 _02178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06360__A2 _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08488__I1 u_arbiter.i_wb_cpu_rdt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06112__A2 _02541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10202__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06240_ u_cpu.rf_ram.memory\[78\]\[2\] _02628_ _02631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07860__A2 _03558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05871__A1 u_cpu.cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06171_ _02585_ _00068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09062__A1 _04294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05122_ _01397_ _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09476__S _04634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07612__A2 _03412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10352__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05623__A1 _01667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05053_ _01544_ _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09930_ _00384_ io_in[4] u_cpu.rf_ram.memory\[57\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09861_ _00315_ io_in[4] u_cpu.rf_ram.memory\[64\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07376__A1 _02832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08812_ _03788_ _03816_ _04246_ _03798_ _04247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_58_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09792_ _00246_ io_in[4] u_cpu.rf_ram.memory\[77\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05926__A2 _02391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09117__A2 _04419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08743_ _03551_ _04199_ _04205_ _01021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05955_ _01403_ _02414_ _02426_ _00010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04906_ _01429_ u_cpu.cpu.state.ibus_cyc _01430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08876__A1 _04292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08674_ u_cpu.cpu.ctrl.o_ibus_adr\[8\] _04155_ _04157_ u_cpu.cpu.ctrl.o_ibus_adr\[9\]
+ _04166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07679__A2 _03454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05886_ u_arbiter.i_wb_cpu_dbus_dat\[5\] _01369_ _02368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07625_ u_cpu.rf_ram.memory\[38\]\[3\] _03422_ _03426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06351__A2 _02695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05785__S1 _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07556_ _03353_ _03382_ _03387_ _00651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__04901__A3 _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06507_ _02746_ _02791_ _02795_ _00194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09718__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06103__A2 _02541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07300__A1 u_cpu.rf_ram.memory\[39\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07487_ _03343_ _03345_ _03346_ _00623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04882__I _01369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09226_ _04476_ _04487_ _04491_ _01218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06438_ _02746_ _02740_ _02747_ _00173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07851__A2 _03558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05862__A1 _02305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09157_ u_cpu.rf_ram.memory\[108\]\[0\] _04449_ _04450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06369_ _02601_ _02637_ _02706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08108_ u_arbiter.i_wb_cpu_dbus_dat\[28\] _03676_ _03721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09868__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07603__A2 _03412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09088_ _04284_ _04409_ _04411_ _01160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08800__A1 _02433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05614__A1 _01398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08039_ _02781_ _03648_ _03675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_1_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10845__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11050_ _11050_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__09356__A2 _04556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07367__A1 _03165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10001_ _00447_ io_in[4] u_cpu.rf_ram.memory\[142\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09108__A2 _04419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06590__A2 _02834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08867__A1 _04286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10903_ _01332_ io_in[4] u_cpu.rf_ram.memory\[98\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06342__A2 _02686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05776__S1 _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10225__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10834_ _01263_ io_in[4] u_cpu.rf_ram.memory\[87\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06049__I _02501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10765_ _01194_ io_in[4] u_cpu.rf_ram.memory\[108\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10696_ _01125_ io_in[4] u_cpu.rf_ram.memory\[102\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10375__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[53\] u_scanchain_local.module_data_in\[52\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[15\] u_scanchain_local.clk u_scanchain_local.module_data_in\[53\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__09044__A1 _04294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09347__A2 _04556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07358__A1 _02602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05128__I _01548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06581__A2 _02834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05740_ _02218_ _02220_ _02222_ _02224_ _01568_ _02225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_76_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05572__B _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08858__A1 _02475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07905__I0 _02587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05671_ u_cpu.rf_ram.memory\[40\]\[6\] u_cpu.rf_ram.memory\[41\]\[6\] u_cpu.rf_ram.memory\[42\]\[6\]
+ u_cpu.rf_ram.memory\[43\]\[6\] _01545_ _01642_ _02157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_36_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07530__A1 _03343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07410_ u_cpu.rf_ram.memory\[133\]\[7\] _03295_ _03303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08390_ u_arbiter.i_wb_cpu_rdt\[27\] u_arbiter.i_wb_cpu_rdt\[11\] _01437_ _03963_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10718__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04895__A2 _01420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07341_ _03264_ _03265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09283__A1 _04480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08086__A2 _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05519__S1 _01620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06097__A1 _02517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07272_ u_cpu.rf_ram.memory\[138\]\[1\] _03225_ _03227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09011_ _02602_ _04197_ _04368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06223_ _02502_ _02614_ _02619_ _00086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10868__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06154_ _02517_ _02563_ _02571_ _00065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05105_ _01397_ _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06085_ _02487_ _02530_ _02532_ _00035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09338__A2 _04546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09913_ _00367_ io_in[4] u_cpu.rf_ram.memory\[5\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05036_ u_arbiter.i_wb_cpu_dbus_adr\[29\] _01457_ _01531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05072__A2 _01414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07349__A1 _03165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09844_ _00298_ io_in[4] u_cpu.rf_ram.memory\[66\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09775_ _00229_ io_in[4] u_cpu.rf_ram.memory\[129\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06987_ _02963_ _03061_ _03066_ _00403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10248__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08726_ _04192_ _04193_ _04194_ _04195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__04877__I _01368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05938_ _02321_ u_cpu.rf_ram.rdata\[3\] _02416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09510__A2 _04654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08657_ _04156_ _04157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05869_ _02309_ _02325_ _02351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06324__A2 _02673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07521__A1 u_cpu.rf_ram.memory\[128\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07608_ _03351_ _03412_ _03416_ _00674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_41_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08588_ _04116_ _00955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_42_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10398__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04886__A2 u_cpu.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07539_ u_cpu.rf_ram.memory\[127\]\[5\] _03372_ _03378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08077__A2 _03683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09690__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10550_ _00982_ io_in[4] u_cpu.rf_ram.memory\[30\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09209_ u_cpu.rf_ram.memory\[84\]\[5\] _04470_ _04481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05835__A1 _02311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09026__A1 _04294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10481_ _00914_ io_in[4] u_cpu.cpu.immdec.imm30_25\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08234__C1 _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07588__A1 _03349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11102_ _11102_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__06260__A1 _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09329__A2 _04546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11033_ _11033_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__08001__A2 _03636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05446__S0 _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06563__A2 _02823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07760__A1 _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05392__B _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09501__A2 _04644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06315__A2 _02673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07512__A1 _03343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10817_ _01246_ io_in[4] u_cpu.rf_ram.memory\[110\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09265__A1 _04480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10748_ _01177_ io_in[4] u_cpu.rf_ram.memory\[107\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07815__A2 _03530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05826__A1 _02309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10679_ _01108_ io_in[4] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08240__A2 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06251__A1 _02517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06910_ _02584_ u_cpu.rf_ram.memory\[5\]\[2\] _03021_ _03024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07890_ _02590_ u_cpu.rf_ram.memory\[8\]\[4\] _03577_ _03582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05437__S0 _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07051__I0 _02581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06841_ u_cpu.rf_ram.memory\[62\]\[3\] _02982_ _02986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07751__A1 u_cpu.rf_ram.memory\[92\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06554__A2 _02821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09560_ _03797_ _03458_ _04683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06772_ _02943_ _02944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08511_ _02768_ _04070_ _04071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05723_ u_cpu.rf_ram.memory\[140\]\[6\] u_cpu.rf_ram.memory\[141\]\[6\] u_cpu.rf_ram.memory\[142\]\[6\]
+ u_cpu.rf_ram.memory\[143\]\[6\] _01680_ _01681_ _02209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09491_ _04468_ _04644_ _04645_ _01329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10540__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06306__A2 _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08700__B1 _04175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08442_ _02433_ _02392_ _03797_ _04011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05514__B1 _01999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05654_ _01570_ _02139_ _02140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05904__I2 u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08373_ _02305_ _03947_ _03948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05585_ u_cpu.rf_ram.memory\[44\]\[5\] u_cpu.rf_ram.memory\[45\]\[5\] u_cpu.rf_ram.memory\[46\]\[5\]
+ u_cpu.rf_ram.memory\[47\]\[5\] _01615_ _01616_ _02072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_51_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10690__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07324_ u_cpu.rf_ram.memory\[49\]\[0\] _03255_ _03256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07806__A2 _03530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09008__A1 _04294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07255_ _03217_ _00520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06206_ _02609_ _00079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05293__A2 _01782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09559__A2 _04674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07186_ _03163_ _03176_ _03179_ _00489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06137_ _02528_ _02561_ _02562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08231__A2 _03778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06068_ u_cpu.rf_ram.memory\[82\]\[7\] _02477_ _02518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07990__A1 _03539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06793__A2 _02955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09906__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05019_ u_cpu.cpu.ctrl.o_ibus_adr\[25\] _01517_ _01518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10070__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09827_ _00281_ io_in[4] u_cpu.rf_ram.memory\[68\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05348__A3 _01837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06545__A2 _02812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09758_ _00212_ io_in[4] u_cpu.rf_ram.memory\[40\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08709_ _04184_ _01008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08298__A2 _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09495__A1 _04474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09689_ _00143_ io_in[4] u_cpu.rf_ram.memory\[41\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05600__S0 _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08028__B _02781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10602_ _01031_ io_in[4] u_cpu.rf_ram.memory\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[41\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05808__A1 _02273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10533_ _00966_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06481__A1 u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10464_ _00897_ io_in[4] u_cpu.rf_ram.memory\[114\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05387__B _01565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10395_ _00828_ io_in[4] u_cpu.rf_ram.memory\[116\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08222__A2 _03742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10413__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07158__I _02486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05036__A2 _01457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09586__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06784__A2 _02944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_scanchain_local.scan_flop\[16\] u_arbiter.i_wb_cpu_rdt\[13\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[10\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
X_11016_ _11016_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_38_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10563__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07733__A1 _02309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08289__A2 _02821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05370_ _01399_ _01859_ _01860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08461__A2 _03786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06472__A1 u_cpu.cpu.state.genblk1.misalign_trap_sync_r vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07040_ u_cpu.rf_ram.memory\[52\]\[4\] _03091_ _03096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05275__A2 _01765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09929__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10093__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09410__A1 _04478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09484__S _04634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08991_ u_cpu.rf_ram.memory\[101\]\[7\] _04349_ _04357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10906__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07972__A1 _03539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06775__A2 _02944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07942_ _03547_ _03606_ _03610_ _00815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07873_ u_cpu.rf_ram.memory\[121\]\[4\] _03568_ _03573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06527__A2 _02801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08772__I0 _02587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09612_ _00066_ io_in[4] u_cpu.rf_ram.memory\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06824_ _02961_ _02972_ _02976_ _00330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09543_ _04673_ _04674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06755_ u_cpu.rf_ram.memory\[65\]\[0\] _02934_ _02935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05706_ _01609_ _02191_ _02192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09474_ _02581_ u_cpu.rf_ram.memory\[0\]\[1\] _04634_ _04636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_70_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06686_ _02896_ _00272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_36_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[64\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08425_ _02392_ _03994_ _03995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05637_ u_cpu.rf_ram.memory\[128\]\[5\] u_cpu.rf_ram.memory\[129\]\[5\] u_cpu.rf_ram.memory\[130\]\[5\]
+ u_cpu.rf_ram.memory\[131\]\[5\] _01687_ _01688_ _02124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09229__A1 u_cpu.rf_ram.memory\[59\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08356_ u_cpu.cpu.immdec.imm24_20\[3\] _03916_ _03933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05568_ _01562_ _02054_ _01582_ _02055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07307_ _03157_ _03245_ _03246_ _00543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08287_ _03816_ _03867_ _03875_ _03876_ _03877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05499_ u_cpu.rf_ram.memory\[36\]\[4\] u_cpu.rf_ram.memory\[37\]\[4\] u_cpu.rf_ram.memory\[38\]\[4\]
+ u_cpu.rf_ram.memory\[39\]\[4\] _01619_ _01620_ _01987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08452__A2 _03797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10436__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07238_ _03161_ _03206_ _03208_ _00512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07169_ _03167_ _03159_ _03168_ _00483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08204__A2 _03802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06215__A1 _02482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07907__S _03586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10180_ _00626_ io_in[4] u_cpu.rf_ram.memory\[22\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10586__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06766__A2 _02934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07715__A1 _03347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06518__A2 _02801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08763__I0 _02599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07191__A2 _03176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09468__A1 _04482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08443__A2 _02305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10516_ _00949_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10929__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10447_ _00880_ io_in[4] u_cpu.rf_ram.memory\[113\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07254__I0 _02581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10378_ _00811_ io_in[4] u_cpu.rf_ram.memory\[112\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07954__A1 _03539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06757__A2 _02934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05965__B1 _01409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05564__C _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06509__A2 _02791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04870_ _01389_ _01391_ _01395_ _01396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_66_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05136__I _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07182__A2 _03176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10309__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06540_ _02742_ _02812_ _02814_ _00208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06168__S _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09601__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08131__A1 _03547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06471_ _02767_ _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08682__A2 _04155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08210_ _03752_ _03800_ _03807_ _03808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__10459__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05496__A2 _01983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05422_ u_cpu.rf_ram.memory\[100\]\[3\] u_cpu.rf_ram.memory\[101\]\[3\] u_cpu.rf_ram.memory\[102\]\[3\]
+ u_cpu.rf_ram.memory\[103\]\[3\] _01577_ _01549_ _01911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_60_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09190_ _04296_ _04459_ _04467_ _01206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08141_ u_arbiter.i_wb_cpu_rdt\[11\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[11\]
+ _01434_ _03741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_53_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05353_ u_cpu.rf_ram.memory\[80\]\[2\] u_cpu.rf_ram.memory\[81\]\[2\] u_cpu.rf_ram.memory\[82\]\[2\]
+ u_cpu.rf_ram.memory\[83\]\[2\] _01590_ _01642_ _01843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09751__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08434__A2 _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08072_ u_arbiter.i_wb_cpu_rdt\[14\] _03653_ _03654_ u_arbiter.i_wb_cpu_dbus_dat\[14\]
+ _03676_ u_arbiter.i_wb_cpu_dbus_dat\[15\] _03698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_05284_ _01684_ _01774_ _01582_ _01775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06996__A2 _03071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07023_ _02963_ _03081_ _03086_ _00419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_127_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06748__A2 _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08974_ _04347_ _01110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07925_ u_cpu.rf_ram.memory\[112\]\[4\] _03596_ _03601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06430__I _02486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07856_ _03549_ _03558_ _03563_ _00776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05046__I _01538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08370__A1 _03831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08370__B2 _03940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06807_ u_cpu.rf_ram.memory\[29\]\[5\] _02955_ _02966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05184__A1 _01636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07787_ u_cpu.rf_ram.memory\[34\]\[1\] _03520_ _03522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04999_ _01445_ _01501_ _01502_ u_arbiter.o_wb_cpu_adr\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09526_ u_cpu.rf_ram.memory\[89\]\[0\] _04664_ _04665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06738_ _02738_ _02924_ _02925_ _00295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__04931__A1 _01445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08122__A1 _02539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09457_ u_cpu.rf_ram.memory\[24\]\[1\] _04625_ _04627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06669_ u_cpu.rf_ram.memory\[75\]\[2\] _02884_ _02887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08408_ _02765_ u_arbiter.i_wb_cpu_rdt\[29\] _03978_ _03979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09388_ _02348_ _04586_ _01429_ _04587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08339_ _03916_ _03917_ _03918_ _03855_ _00904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_137_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05239__A2 _01725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10301_ _00734_ io_in[4] u_cpu.rf_ram.memory\[92\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06987__A2 _03061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10232_ _00672_ io_in[4] u_cpu.rf_ram.memory\[123\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07936__A1 _03539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06739__A2 _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05665__B _01564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10163_ _00609_ io_in[4] u_cpu.rf_ram.memory\[130\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10094_ _00540_ io_in[4] u_cpu.rf_ram.memory\[39\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_scanchain_local.scan_flop\[9\] u_arbiter.i_wb_cpu_rdt\[6\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[3\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_48_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09624__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08361__A1 _03755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05270__S1 _01668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10601__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10996_ _10996_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_16_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09774__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08664__A2 _04155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10751__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08416__A2 _03751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07475__I0 _02590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06978__A2 _03061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05089__S1 _01580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05971_ _02436_ _01431_ u_arbiter.o_wb_cpu_we vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10131__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07710_ _02475_ _02638_ _03474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04922_ u_arbiter.i_wb_cpu_dbus_adr\[2\] _01443_ _01444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08690_ _04174_ _00999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_39_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08352__A1 _03890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07641_ u_cpu.rf_ram.memory\[37\]\[2\] _03432_ _03435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04853_ _01371_ _01378_ _01379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_26_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06902__A2 _03012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10281__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07572_ _03351_ _03392_ _03396_ _00658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05261__S1 _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08104__A1 u_arbiter.i_wb_cpu_rdt\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09311_ _04472_ _04536_ _04538_ _01256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06523_ _02744_ _02801_ _02804_ _00201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05469__A2 _01956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09242_ _02587_ u_cpu.rf_ram.memory\[10\]\[3\] _04496_ _04500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06666__A1 _02738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06454_ _02581_ u_cpu.rf_ram.memory\[4\]\[1\] _02756_ _02758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05405_ _01601_ _01893_ _01605_ _01894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09173_ _02524_ _02626_ _04458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06385_ _02512_ _02708_ _02715_ _00152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08407__A2 u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08124_ u_cpu.rf_ram.memory\[113\]\[0\] _03731_ _03732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06418__A1 _02502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05336_ u_cpu.rf_ram.memory\[96\]\[2\] u_cpu.rf_ram.memory\[97\]\[2\] u_cpu.rf_ram.memory\[98\]\[2\]
+ u_cpu.rf_ram.memory\[99\]\[2\] _01602_ _01579_ _01826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_108_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06425__I _02481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09080__A2 _04399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06969__A2 _03051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08055_ u_arbiter.i_wb_cpu_rdt\[8\] _03669_ _03678_ u_arbiter.i_wb_cpu_dbus_dat\[8\]
+ _03687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07091__A1 _02961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05267_ u_cpu.rf_ram.memory\[84\]\[1\] u_cpu.rf_ram.memory\[85\]\[1\] u_cpu.rf_ram.memory\[86\]\[1\]
+ u_cpu.rf_ram.memory\[87\]\[1\] _01555_ _01652_ _01758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_134_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07006_ u_cpu.rf_ram.memory\[54\]\[5\] _03071_ _03077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05198_ _01399_ _01689_ _01690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07918__A1 _03539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09647__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07394__A2 _02832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06160__I _02576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08957_ u_arbiter.i_wb_cpu_rdt\[23\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[7\]
+ _04331_ _04339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_u_scanchain_local.scan_flop\[32\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07908_ _03591_ _00800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10624__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08888_ _04284_ _04299_ _04301_ _01070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05157__A1 _01645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07839_ _02511_ _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09797__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08894__A2 _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10850_ _01279_ io_in[4] u_cpu.cpu.genblk3.csr.mcause3_0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[47\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09509_ _04468_ _04654_ _04655_ _01337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_112_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10781_ _01210_ io_in[4] u_cpu.rf_ram.memory\[84\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10774__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08646__A2 _04145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10004__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08751__S _04208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05880__A2 u_cpu.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09071__A2 _04399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07082__A1 _02625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10154__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08957__I0 u_arbiter.i_wb_cpu_rdt\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10215_ _00661_ io_in[4] u_cpu.rf_ram.memory\[125\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07385__A2 _03285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10146_ _00592_ io_in[4] u_cpu.rf_ram.memory\[132\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05396__A1 _01542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10077_ _00523_ io_in[4] u_cpu.rf_ram.memory\[14\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08334__A1 _02436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05148__A1 _01601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08885__A2 _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06896__A1 _02961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10979_ _10979_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_16_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06648__A1 _02738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05320__A1 _01609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06170_ _02584_ u_cpu.rf_ram.memory\[1\]\[2\] _02578_ _02585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05289__C _01404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09062__A2 _04389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05121_ _01609_ _01612_ _01613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05052_ _01543_ _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06820__A1 _02957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05623__A2 _02109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09860_ _00314_ io_in[4] u_cpu.rf_ram.memory\[64\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10647__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07376__A2 _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08811_ u_cpu.cpu.immdec.imm11_7\[1\] u_cpu.cpu.immdec.imm11_7\[2\] _04236_ _04246_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_98_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09791_ _00245_ io_in[4] u_cpu.rf_ram.memory\[77\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05387__A1 _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05926__A3 _02406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08742_ u_cpu.rf_ram.memory\[109\]\[5\] _04199_ _04205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05954_ u_cpu.rf_ram_if.rdata0\[3\] _01403_ _02426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08325__A1 _03831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07128__A2 _03139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_04905_ _01428_ _01429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_54_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08673_ _04165_ _00991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_54_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05139__A1 _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10797__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05885_ _01373_ _01370_ _02367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_54_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08876__A2 _04282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07624_ _03349_ _03422_ _03425_ _00681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06887__A1 _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07555_ u_cpu.rf_ram.memory\[126\]\[4\] _03382_ _03387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08089__B1 _03654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10027__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04901__A4 _01426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06506_ u_cpu.rf_ram.memory\[16\]\[3\] _02791_ _02795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07486_ u_cpu.rf_ram.memory\[22\]\[0\] _03345_ _03346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07300__A2 _03235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09225_ u_cpu.rf_ram.memory\[59\]\[3\] _04487_ _04491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06437_ u_cpu.rf_ram.memory\[50\]\[3\] _02740_ _02747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05311__A1 _01589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09156_ _04448_ _04449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05862__A2 _02344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06368_ _02517_ _02697_ _02705_ _00145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09053__A2 _04389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10177__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08107_ _03717_ _03678_ _03720_ _00870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05319_ u_cpu.rf_ram.memory\[40\]\[2\] u_cpu.rf_ram.memory\[41\]\[2\] u_cpu.rf_ram.memory\[42\]\[2\]
+ u_cpu.rf_ram.memory\[43\]\[2\] _01610_ _01611_ _01809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09087_ u_cpu.rf_ram.memory\[105\]\[1\] _04409_ _04411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06299_ _02492_ _02662_ _02665_ _00116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08800__A2 _02453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08038_ _02774_ _03673_ _03674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06811__A1 _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05170__S0 _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07367__A2 _03275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10000_ _00007_ io_in[4] u_cpu.rf_ram.rdata\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05378__A1 _01858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09989_ _00443_ io_in[4] u_cpu.rf_ram.memory\[15\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08316__A1 _03785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06178__I0 _02590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08867__A2 _04282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10902_ _01331_ io_in[4] u_cpu.rf_ram.memory\[98\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06878__A1 _02961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10833_ _01262_ io_in[4] u_cpu.rf_ram.memory\[111\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05550__A1 _01399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10764_ _01193_ io_in[4] u_cpu.rf_ram.memory\[108\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09292__A2 _04526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05302__A1 _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10695_ _01124_ io_in[4] u_cpu.rf_ram.memory\[102\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09812__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09044__A2 _04379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[46\] u_scanchain_local.module_data_in\[45\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[8\] u_scanchain_local.clk u_scanchain_local.module_data_in\[46\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_126_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06802__A1 _02961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05161__S0 _01623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09962__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07358__A2 _02832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08555__A1 _03549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10129_ _00575_ io_in[4] u_cpu.rf_ram.memory\[134\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08858__A2 _02625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06869__A1 _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05670_ _02149_ _02151_ _02153_ _02155_ _01607_ _02156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_91_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05144__I _01397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07530__A2 _03372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05541__A1 _01636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07340_ _02810_ _02832_ _03264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06176__S _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09283__A2 _04516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07294__A1 u_cpu.rf_ram.memory\[39\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07271_ _03157_ _03225_ _03226_ _00527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06097__A2 _02530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09010_ _04296_ _04359_ _04367_ _01126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06222_ u_cpu.rf_ram.memory\[80\]\[4\] _02614_ _02619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09035__A2 _04379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06153_ u_cpu.rf_ram.memory\[20\]\[7\] _02563_ _02571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07597__A2 _03402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05104_ _01594_ _01595_ _01564_ _01596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_132_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06084_ u_cpu.rf_ram.memory\[21\]\[1\] _02530_ _02532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05035_ u_cpu.cpu.ctrl.o_ibus_adr\[29\] _01529_ _01530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09912_ _00366_ io_in[4] u_cpu.rf_ram.memory\[19\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07349__A2 _03265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09843_ _00297_ io_in[4] u_cpu.rf_ram.memory\[66\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06986_ u_cpu.rf_ram.memory\[55\]\[4\] _03061_ _03066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09774_ _00228_ io_in[4] u_cpu.rf_ram.memory\[129\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08725_ _02324_ _02356_ _04192_ _04194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05937_ _02320_ _02414_ _02415_ _00016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05780__A1 _01589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08849__A2 _04271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08656_ _01428_ _02449_ _04156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08566__S _02445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05868_ _02349_ _02350_ u_cpu.cpu.o_wdata1 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05054__I _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07521__A2 _03362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07607_ u_cpu.rf_ram.memory\[123\]\[3\] _03412_ _03416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05532__A1 _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08587_ u_arbiter.i_wb_cpu_dbus_adr\[14\] u_arbiter.i_wb_cpu_dbus_adr\[13\] _04115_
+ _04116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05799_ _01667_ _02283_ _02284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07538_ _03353_ _03372_ _03377_ _00643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09274__A2 _04516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09835__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06088__A2 _02530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07285__A1 _03173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07469_ _02581_ u_cpu.rf_ram.memory\[12\]\[1\] _03334_ _03336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09208_ _02506_ _04480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10812__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10480_ _00913_ io_in[4] u_cpu.cpu.immdec.imm30_25\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09026__A2 _04369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05391__S0 _01578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09139_ u_cpu.rf_ram.memory\[83\]\[0\] _04439_ _04440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07037__A1 _02959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08234__B1 _03818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09985__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08234__C2 _03802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09196__I _02486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07588__A2 _03402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08785__A1 _03539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05599__A1 _01636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11101_ _11101_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_78_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06260__A2 _02641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[2\]_D u_arbiter.i_wb_cpu_ack vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08537__A1 _03549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11032_ _11032_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_2_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05446__S1 _01668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07760__A2 _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05771__A1 _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07899__I0 _02573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07512__A2 _03362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10342__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05523__B2 _02010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10816_ _01245_ io_in[4] u_cpu.rf_ram.memory\[110\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09265__A2 _04506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08473__B1 _04035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10747_ _01176_ io_in[4] u_cpu.rf_ram.memory\[107\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10492__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09017__A2 _04369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10678_ _01107_ io_in[4] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05382__S0 _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08225__B1 _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07579__A2 _03392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06251__A2 _02628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09708__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06840_ _02959_ _02982_ _02985_ _00337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07200__A1 _03157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05437__S1 _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07751__A2 _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06771_ _02612_ _02626_ _02943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05762__A1 _01397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08510_ _01437_ u_arbiter.i_wb_cpu_rdt\[19\] _03782_ _04069_ _04070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05722_ _01399_ _02207_ _02208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09490_ u_cpu.rf_ram.memory\[98\]\[0\] _04644_ _04645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09858__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08441_ _03744_ _03816_ _04009_ _03876_ _04010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_1_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05653_ u_cpu.rf_ram.memory\[20\]\[6\] u_cpu.rf_ram.memory\[21\]\[6\] u_cpu.rf_ram.memory\[22\]\[6\]
+ u_cpu.rf_ram.memory\[23\]\[6\] _01572_ _01574_ _02139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05904__I3 u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08372_ _02436_ _02313_ _02434_ _03947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10835__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05584_ _01609_ _02070_ _02071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09256__A2 _04506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07323_ _03254_ _03255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07254_ _02581_ u_cpu.rf_ram.memory\[14\]\[1\] _03215_ _03217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09008__A2 _04359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05373__S0 _01687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06205_ _02593_ u_cpu.rf_ram.memory\[7\]\[5\] _02603_ _02609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07019__A1 _02959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07185_ u_cpu.rf_ram.memory\[73\]\[2\] _03176_ _03179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06136_ _02523_ _02560_ _02561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06433__I _02491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05125__S0 _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06242__A2 _02628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06067_ _02516_ _02517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10215__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05049__I _01540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07990__A2 _03636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05018_ u_cpu.cpu.ctrl.o_ibus_adr\[24\] _01513_ _01517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09192__A1 _02475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05493__B _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09826_ _00280_ io_in[4] u_cpu.rf_ram.memory\[68\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10365__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09757_ _00211_ io_in[4] u_cpu.rf_ram.memory\[40\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05753__A1 _01540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06969_ _02963_ _03051_ _03056_ _00395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08708_ u_cpu.cpu.ctrl.o_ibus_adr\[24\] _04173_ _04175_ u_cpu.cpu.ctrl.o_ibus_adr\[25\]
+ _04184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09688_ _00142_ io_in[4] u_cpu.rf_ram.memory\[41\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09495__A2 _04644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05505__A1 _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08639_ _03539_ _04145_ _04146_ _00976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_54_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05600__S1 _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10601_ _01030_ io_in[4] u_cpu.rf_ram.memory\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10532_ _00965_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05364__S0 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10463_ _00896_ io_in[4] u_cpu.rf_ram.memory\[114\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10394_ _00827_ io_in[4] u_cpu.rf_ram.memory\[115\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07430__A1 _02682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07981__A2 _03626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10708__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05992__A1 _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11015_ _11015_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_89_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05744__A1 _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10858__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08694__B1 _04175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06454__S _02756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05355__S0 _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10238__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05107__S0 _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09410__A2 _04595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06224__A2 _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07421__A1 _03165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08990_ _04294_ _04349_ _04356_ _01117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07972__A2 _03626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07941_ u_cpu.rf_ram.memory\[122\]\[3\] _03606_ _03610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10388__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05983__A1 u_cpu.cpu.genblk3.csr.o_new_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07872_ _03547_ _03568_ _03572_ _00783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07724__A2 _03475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08921__A1 u_arbiter.i_wb_cpu_ack vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09680__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09611_ _00065_ io_in[4] u_cpu.rf_ram.memory\[20\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06823_ u_cpu.rf_ram.memory\[63\]\[3\] _02972_ _02976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05735__A1 _01398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09542_ _02528_ _02602_ _04673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06754_ _02933_ _02934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05705_ u_cpu.rf_ram.memory\[80\]\[6\] u_cpu.rf_ram.memory\[81\]\[6\] u_cpu.rf_ram.memory\[82\]\[6\]
+ u_cpu.rf_ram.memory\[83\]\[6\] _01590_ _01591_ _02191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_36_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06685_ _02581_ u_cpu.rf_ram.memory\[6\]\[1\] _02894_ _02896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09473_ _04635_ _01321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08424_ _01372_ _02313_ u_cpu.cpu.decode.opcode\[1\] _03994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05636_ _01684_ _02122_ _01582_ _02123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_u_scanchain_local.scan_flop\[26\]_D u_arbiter.i_wb_cpu_rdt\[23\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05594__S0 _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09229__A2 _04487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08355_ u_cpu.cpu.immdec.imm24_20\[4\] _02768_ _03932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05567_ u_cpu.rf_ram.memory\[16\]\[5\] u_cpu.rf_ram.memory\[17\]\[5\] u_cpu.rf_ram.memory\[18\]\[5\]
+ u_cpu.rf_ram.memory\[19\]\[5\] _01578_ _01580_ _02054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08988__A1 _04292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07306_ u_cpu.rf_ram.memory\[137\]\[0\] _03245_ _03246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08286_ _03796_ _03782_ _03876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_109_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05498_ _01397_ _01985_ _01605_ _01986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_109_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07237_ u_cpu.rf_ram.memory\[143\]\[1\] _03206_ _03208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07660__A1 _03349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07168_ u_cpu.rf_ram.memory\[72\]\[4\] _03159_ _03168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09401__A2 _04595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06215__A2 _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07412__A1 _02561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06119_ u_cpu.rf_ram.memory\[18\]\[0\] _02551_ _02552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07099_ _02969_ _03119_ _03127_ _00454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07963__A2 _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05974__A1 _02309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07715__A2 _03475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08912__A1 _04290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09809_ _00263_ io_in[4] u_cpu.rf_ram.memory\[75\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05726__A1 _01399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09468__A2 _04625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08676__B1 _04157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05670__C _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[17\]_D u_arbiter.i_wb_cpu_rdt\[14\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05585__S0 _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10515_ _00948_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10446_ _00879_ io_in[4] u_cpu.rf_ram.memory\[113\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10530__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07403__A1 _03165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10377_ _00810_ io_in[4] u_cpu.rf_ram.memory\[112\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07954__A2 _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05965__A1 _02332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05965__B2 _02361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08203__I0 u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10680__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07706__A2 _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05717__A1 _01553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09459__A2 _04625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04940__A2 _01457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08131__A2 _03731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06470_ _02765_ u_arbiter.i_wb_cpu_ibus_adr\[1\] _02766_ _02767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_61_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06142__A1 _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05576__S0 _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05421_ _01594_ _01909_ _01416_ _01910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_53_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10060__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08140_ _02768_ _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05352_ _01645_ _01841_ _01648_ _01842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_105_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06184__S _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07642__A1 _03349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08071_ _03696_ _03697_ _00857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05283_ u_cpu.rf_ram.memory\[140\]\[1\] u_cpu.rf_ram.memory\[141\]\[1\] u_cpu.rf_ram.memory\[142\]\[1\]
+ u_cpu.rf_ram.memory\[143\]\[1\] _01680_ _01681_ _01774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_128_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07022_ u_cpu.rf_ram.memory\[53\]\[4\] _03081_ _03086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06912__S _03021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09395__A1 u_cpu.cpu.ctrl.i_iscomp vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07945__A2 _03606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08973_ u_arbiter.i_wb_cpu_rdt\[31\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\]
+ _04331_ _04347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07924_ _03547_ _03596_ _03600_ _00807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[31\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07855_ u_cpu.rf_ram.memory\[118\]\[4\] _03558_ _03563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05708__A1 _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08370__A2 _03773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06806_ _02506_ _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07786_ _03343_ _03520_ _03521_ _00748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06381__A1 _02502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04998_ u_arbiter.i_wb_cpu_dbus_adr\[20\] _01457_ _01502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09525_ _04663_ _04664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08658__B1 _04157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06737_ u_cpu.rf_ram.memory\[66\]\[0\] _02924_ _02925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08122__A2 _02821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10403__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08574__S _02445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09456_ _04468_ _04625_ _04626_ _01313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06668_ _02742_ _02884_ _02886_ _00264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05567__S0 _01578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05062__I _01553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09576__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05619_ u_cpu.rf_ram.memory\[84\]\[5\] u_cpu.rf_ram.memory\[85\]\[5\] u_cpu.rf_ram.memory\[86\]\[5\]
+ u_cpu.rf_ram.memory\[87\]\[5\] _01555_ _01652_ _02106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_12_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08407_ _01437_ u_arbiter.i_wb_cpu_rdt\[13\] _03978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__07881__A1 _02577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09387_ _02339_ _03454_ _04585_ _04586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06599_ u_cpu.rf_ram.memory\[139\]\[3\] _02844_ _02848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08338_ u_cpu.cpu.immdec.imm24_20\[0\] _03916_ _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05319__S0 _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10553__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08269_ _03767_ _03768_ _03860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_125_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10300_ _00733_ io_in[4] u_cpu.rf_ram.memory\[92\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04998__A2 _01457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10231_ _00671_ io_in[4] u_cpu.rf_ram.memory\[123\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08189__A2 _03788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09386__A1 u_cpu.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07936__A2 _03606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10162_ _00608_ io_in[4] u_cpu.rf_ram.memory\[130\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05947__A1 _02321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08041__C _03676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10093_ _00539_ io_in[4] u_cpu.rf_ram.memory\[39\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08749__S _04208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08361__A2 _03757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04922__A2 _01443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10995_ _10995_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__09919__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08113__A2 _03718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10083__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06124__A1 _02492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05558__S0 _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07872__A1 _03547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06675__A2 _02884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07624__A1 _03349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09377__A1 _01381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10429_ _00862_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07927__A2 _03596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[54\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05938__A1 _02321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05970_ _02306_ _02436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_97_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04921_ _01442_ _01443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08352__A2 _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07640_ _03347_ _03432_ _03434_ _00688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10426__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04852_ _01372_ _01374_ _01378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07571_ u_cpu.rf_ram.memory\[125\]\[3\] _03392_ _03396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09599__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09301__A1 _04480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08104__A2 _03653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09310_ u_cpu.rf_ram.memory\[111\]\[1\] _04536_ _04538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06522_ u_cpu.rf_ram.memory\[17\]\[2\] _02801_ _02804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05549__S0 _01687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10576__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09241_ _04499_ _01225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06453_ _02757_ _00178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07863__A1 _02695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06666__A2 _02884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06910__I0 _02584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05404_ u_cpu.rf_ram.memory\[56\]\[3\] u_cpu.rf_ram.memory\[57\]\[3\] u_cpu.rf_ram.memory\[58\]\[3\]
+ u_cpu.rf_ram.memory\[59\]\[3\] _01602_ _01579_ _01893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09172_ _04296_ _04449_ _04457_ _01198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06384_ u_cpu.rf_ram.memory\[43\]\[6\] _02708_ _02715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08123_ _03730_ _03731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06418__A2 _02729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05335_ _01636_ _01824_ _01825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08054_ u_arbiter.i_wb_cpu_dbus_dat\[9\] _03683_ _03686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05266_ _01609_ _01756_ _01757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07091__A2 _03119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05721__S0 _01687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09368__A1 _02341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07005_ _02963_ _03071_ _03076_ _00411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05766__B _01626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08415__I0 u_arbiter.i_wb_cpu_rdt\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05197_ u_cpu.rf_ram.memory\[128\]\[0\] u_cpu.rf_ram.memory\[129\]\[0\] u_cpu.rf_ram.memory\[130\]\[0\]
+ u_cpu.rf_ram.memory\[131\]\[0\] _01687_ _01688_ _01689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_131_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07918__A2 _03596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05929__A1 _01374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05485__C _01426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08956_ _04338_ _01101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05057__I _01548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07473__S _03334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07907_ _02590_ u_cpu.rf_ram.memory\[11\]\[4\] _03586_ _03591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_57_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08887_ u_cpu.rf_ram.memory\[95\]\[1\] _04299_ _04301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04896__I _01421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07838_ _03551_ _03541_ _03552_ _00769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05157__A2 _01647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06354__A1 _02482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07769_ u_cpu.rf_ram.memory\[35\]\[1\] _03510_ _03512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10919__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09508_ u_cpu.rf_ram.memory\[100\]\[0\] _04654_ _04655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06106__A1 _02492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10780_ _01209_ io_in[4] u_cpu.rf_ram.memory\[84\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07854__A1 _03547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06657__A2 _02874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09439_ u_cpu.rf_ram.memory\[25\]\[1\] _04615_ _04617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09199__I _02491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07606__A1 _03349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06409__A2 _02729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05880__A3 _01385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07082__A2 _02832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05712__S0 _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05093__A1 _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09359__A1 _04484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10214_ _00660_ io_in[4] u_cpu.rf_ram.memory\[125\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10145_ _00591_ io_in[4] u_cpu.rf_ram.memory\[132\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10449__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05235__I3 u_cpu.rf_ram.memory\[39\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05396__A2 _01884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10076_ _00522_ io_in[4] u_cpu.rf_ram.memory\[14\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09531__A1 _04474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08334__A2 _02313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09741__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05148__A2 _01639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06345__A1 _02507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05779__S0 _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10599__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06896__A2 _03012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10978_ _10978_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_15_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07145__I0 _02590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09891__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07845__A1 _02821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06648__A2 _02874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05320__A2 _01809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05120_ u_cpu.rf_ram.memory\[40\]\[0\] u_cpu.rf_ram.memory\[41\]\[0\] u_cpu.rf_ram.memory\[42\]\[0\]
+ u_cpu.rf_ram.memory\[43\]\[0\] _01610_ _01611_ _01612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_129_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06462__S _02756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08270__A1 _03768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05703__S0 _01646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05084__A1 _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05051_ u_cpu.raddr\[0\] _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05586__B _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06820__A2 _02972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08022__A1 u_arbiter.i_wb_cpu_rdt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08810_ _03740_ _04242_ _04244_ _04245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09790_ _00244_ io_in[4] u_cpu.rf_ram.memory\[77\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06584__A1 _02748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08741_ _03549_ _04199_ _04204_ _01020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05953_ _01403_ _02412_ _02425_ _00009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08325__A2 _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04904_ io_in[1] _01428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08672_ u_cpu.cpu.ctrl.o_ibus_adr\[7\] _04155_ _04157_ u_cpu.cpu.ctrl.o_ibus_adr\[8\]
+ _04165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05884_ _02305_ _02362_ _02365_ _02366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_66_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05139__A2 _01569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07623_ u_cpu.rf_ram.memory\[38\]\[2\] _03422_ _03425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06887__A2 _02682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08089__A1 u_arbiter.i_wb_cpu_rdt\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07554_ _03351_ _03382_ _03386_ _00650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06505_ _02744_ _02791_ _02794_ _00193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06639__A2 _02864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07485_ _03344_ _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09224_ _04474_ _04487_ _04490_ _01217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06436__I _02496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06436_ _02496_ _02746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05311__A2 _01800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09155_ _02671_ _04197_ _04448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06367_ u_cpu.rf_ram.memory\[41\]\[7\] _02697_ _02705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08106_ u_arbiter.i_wb_cpu_rdt\[26\] _02781_ _03718_ u_arbiter.i_wb_cpu_dbus_dat\[27\]
+ _03720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__09614__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05318_ _01801_ _01803_ _01805_ _01807_ _01607_ _01808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_107_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08261__A1 _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09086_ _04280_ _04409_ _04410_ _01159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06298_ u_cpu.rf_ram.memory\[45\]\[2\] _02662_ _02665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05249_ _01601_ _01739_ _01626_ _01740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08037_ u_arbiter.i_wb_cpu_dbus_dat\[4\] _02775_ _03673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06811__A2 _02955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05170__S1 _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09764__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09988_ _00442_ io_in[4] u_cpu.rf_ram.memory\[15\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05378__A2 _01867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08939_ _04294_ _04322_ _04329_ _01093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10741__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09513__A1 _04474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08316__A2 _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10901_ _01330_ io_in[4] u_cpu.rf_ram.memory\[98\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06878__A2 _03002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10832_ _01261_ io_in[4] u_cpu.rf_ram.memory\[111\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10891__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10763_ _01192_ io_in[4] u_cpu.rf_ram.memory\[108\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10694_ _01123_ io_in[4] u_cpu.rf_ram.memory\[102\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10121__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08252__A1 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06802__A2 _02955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_scanchain_local.scan_flop\[39\] u_scanchain_local.module_data_in\[38\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[1\] u_scanchain_local.clk u_scanchain_local.module_data_in\[39\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__10271__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05161__S1 _01652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08004__A1 _03555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08555__A2 _04094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06566__A1 u_cpu.rf_ram.memory\[119\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08510__B _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10128_ _00574_ io_in[4] u_cpu.rf_ram.memory\[135\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10059_ _00505_ io_in[4] u_cpu.rf_ram.memory\[70\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06318__A1 _02492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06869__A2 _02684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07818__A1 _03359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07270_ u_cpu.rf_ram.memory\[138\]\[0\] _03225_ _03226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09637__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07294__A2 _03235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05160__I _01547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06221_ _02497_ _02614_ _02618_ _00085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_u_scanchain_local.scan_flop\[31\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10614__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06152_ _02512_ _02563_ _02570_ _00064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08243__A1 _03742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07046__A2 _03091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05103_ u_cpu.rf_ram.memory\[48\]\[0\] u_cpu.rf_ram.memory\[49\]\[0\] u_cpu.rf_ram.memory\[50\]\[0\]
+ u_cpu.rf_ram.memory\[51\]\[0\] _01544_ _01548_ _01595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09787__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08794__A2 _04227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06083_ _02482_ _02530_ _02531_ _00034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_u_scanchain_local.scan_flop\[46\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05034_ u_cpu.cpu.ctrl.o_ibus_adr\[28\] u_cpu.cpu.ctrl.o_ibus_adr\[27\] _01523_ _01529_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09911_ _00365_ io_in[4] u_cpu.rf_ram.memory\[19\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06920__S _03021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10764__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08546__A2 _04094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09842_ _00296_ io_in[4] u_cpu.rf_ram.memory\[66\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_101_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06557__A1 _02738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08420__B _03906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09773_ _00227_ io_in[4] u_cpu.rf_ram.memory\[129\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06985_ _02961_ _03061_ _03065_ _00402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08724_ _02381_ _02406_ u_cpu.cpu.ctrl.i_jump _04193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06309__A1 _02517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05936_ _02320_ u_cpu.rf_ram_if.rdata1\[2\] _02415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05780__A2 _02264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08655_ _04154_ _04155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_15_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05867_ u_arbiter.i_wb_cpu_ibus_adr\[0\] _01386_ _02350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07606_ _03349_ _03412_ _03415_ _00673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08586_ _02372_ _04115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05532__A2 _02019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05798_ u_cpu.rf_ram.memory\[64\]\[7\] u_cpu.rf_ram.memory\[65\]\[7\] u_cpu.rf_ram.memory\[66\]\[7\]
+ u_cpu.rf_ram.memory\[67\]\[7\] _01571_ _01668_ _02283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10144__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07537_ u_cpu.rf_ram.memory\[127\]\[4\] _03372_ _03377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08582__S _02445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07468_ _03335_ _00615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07285__A2 _03225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05070__I _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09207_ _04478_ _04470_ _04479_ _01211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06419_ u_cpu.rf_ram.memory\[47\]\[5\] _02729_ _02735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08609__I0 u_arbiter.i_wb_cpu_dbus_adr\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10294__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07399_ _03161_ _03295_ _03297_ _00584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05391__S1 _01580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09138_ _04438_ _04439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08234__A1 _03763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07037__A2 _03091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08785__A2 _04227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09069_ u_cpu.rf_ram.memory\[79\]\[1\] _04399_ _04401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05599__A2 _02085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06796__A1 _02957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11100_ _11100_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_118_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08537__A2 _04084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11031_ _11031_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__06548__A1 _02750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05220__A1 _01542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08757__S _04208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05771__A2 _02255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06720__A1 _02738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10815_ _01244_ io_in[4] u_cpu.rf_ram.memory\[110\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10637__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10746_ _01175_ io_in[4] u_cpu.rf_ram.memory\[107\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08473__A1 _01390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07276__A2 _03225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10677_ _01106_ io_in[4] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05382__S1 _01557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08225__A1 _03754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07028__A2 _03081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08225__B2 _03759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10787__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08528__A2 _04084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10017__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08240__B _03834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07200__A2 _03186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05211__A1 _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06770_ _02754_ _02934_ _02942_ _00310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05762__A2 _02246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10167__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05721_ u_cpu.rf_ram.memory\[136\]\[6\] u_cpu.rf_ram.memory\[137\]\[6\] u_cpu.rf_ram.memory\[138\]\[6\]
+ u_cpu.rf_ram.memory\[139\]\[6\] _01687_ _01681_ _02207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_91_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08440_ _04007_ _04008_ _04009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08700__A2 _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05652_ _02131_ _02133_ _02135_ _02137_ _01568_ _02138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_51_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05583_ u_cpu.rf_ram.memory\[40\]\[5\] u_cpu.rf_ram.memory\[41\]\[5\] u_cpu.rf_ram.memory\[42\]\[5\]
+ u_cpu.rf_ram.memory\[43\]\[5\] _01545_ _01642_ _02070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08371_ _03876_ _03945_ _03946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_51_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07322_ _02539_ _02684_ _03254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05104__B _01564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08464__A1 _04024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07253_ _03216_ _00519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05373__S1 _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06204_ _02608_ _00078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08216__A1 _03773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07019__A2 _03081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07184_ _03161_ _03176_ _03178_ _00488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05758__C _01425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06135_ _01668_ _02466_ _02560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_117_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05125__S1 _01616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06778__A1 _02744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06066_ _02515_ _02516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05017_ _01445_ _01515_ _01516_ u_arbiter.o_wb_cpu_adr\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_63_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09192__A2 _02561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09825_ _00279_ io_in[4] u_cpu.rf_ram.memory\[68\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05202__A1 _01679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09756_ _00210_ io_in[4] u_cpu.rf_ram.memory\[40\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06968_ u_cpu.rf_ram.memory\[56\]\[4\] _03051_ _03056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05065__I _01548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05753__A2 _02237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07481__S _03334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09802__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08707_ _04183_ _01007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05919_ u_cpu.cpu.decode.opcode\[1\] _02313_ _02314_ _02400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09687_ _00141_ io_in[4] u_cpu.rf_ram.memory\[41\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06899_ u_cpu.rf_ram.memory\[19\]\[5\] _03012_ _03018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08638_ u_cpu.rf_ram.memory\[30\]\[0\] _04145_ _04146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05505__A2 _01964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06702__A1 _02738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08569_ _04106_ _00946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09952__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10600_ _01029_ io_in[4] u_cpu.rf_ram.memory\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10531_ _00964_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08325__B _03791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05364__S1 _01549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08207__A1 u_cpu.cpu.decode.opcode\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10462_ _00895_ io_in[4] u_cpu.rf_ram.memory\[114\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10393_ _00826_ io_in[4] u_cpu.rf_ram.memory\[115\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07430__A2 _02832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05992__A2 _02313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11014_ _11014_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__09183__A2 _04459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07194__A1 _03171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08391__B1 _03963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08930__A2 _04322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[5\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07249__A2 _03206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08997__A2 _04359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10729_ _01158_ io_in[4] u_cpu.rf_ram.memory\[79\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05859__B _02338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05355__S1 _01652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09246__I0 _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05680__A1 _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05107__S1 _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07421__A2 _03305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05432__A1 _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07940_ _03545_ _03606_ _03609_ _00814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05983__A2 u_cpu.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09825__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07871_ u_cpu.rf_ram.memory\[121\]\[3\] _03568_ _03572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09610_ _00064_ io_in[4] u_cpu.rf_ram.memory\[20\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06822_ _02959_ _02972_ _02975_ _00329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10802__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09541_ _04484_ _04664_ _04672_ _01352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06753_ _02539_ _02626_ _02933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09975__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05704_ _01645_ _02189_ _01648_ _02190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_110_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09472_ _02573_ u_cpu.rf_ram.memory\[0\]\[0\] _04634_ _04635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06684_ _02895_ _00271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_58_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08423_ u_cpu.cpu.immdec.imm19_12_20\[0\] _03993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05635_ u_cpu.rf_ram.memory\[140\]\[5\] u_cpu.rf_ram.memory\[141\]\[5\] u_cpu.rf_ram.memory\[142\]\[5\]
+ u_cpu.rf_ram.memory\[143\]\[5\] _01680_ _01681_ _02122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_12_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10952__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05594__S1 _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08354_ _03782_ _03923_ _03930_ _03797_ _03931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__08437__A1 _03999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05566_ _01570_ _02052_ _02053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07305_ _03244_ _03245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08988__A2 _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05497_ u_cpu.rf_ram.memory\[44\]\[4\] u_cpu.rf_ram.memory\[45\]\[4\] u_cpu.rf_ram.memory\[46\]\[4\]
+ u_cpu.rf_ram.memory\[47\]\[4\] _01615_ _01616_ _01985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08285_ _03851_ _03872_ _03873_ _03874_ _03875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06999__A1 _02957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07236_ _03157_ _03206_ _03207_ _00511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07660__A2 _03442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07167_ _02501_ _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06118_ _02550_ _02551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07412__A2 _02832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10332__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07098_ u_cpu.rf_ram.memory\[142\]\[7\] _03119_ _03127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05423__A1 _01636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06049_ _02501_ _02502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09165__A2 _04449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08912__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09808_ _00262_ io_in[4] u_cpu.rf_ram.memory\[76\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10482__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09739_ _00193_ io_in[4] u_cpu.rf_ram.memory\[16\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06151__A2 _02563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05585__S1 _01616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08428__A1 _03991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09476__I0 _02584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08979__A2 _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07100__A1 _02660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10514_ _00947_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08770__S _04217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07651__A2 _03432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10445_ _00878_ io_in[4] u_cpu.rf_ram.memory\[113\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09848__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07403__A2 _03295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10376_ _00809_ io_in[4] u_cpu.rf_ram.memory\[112\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05414__A1 _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06462__I0 _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[21\] u_arbiter.i_wb_cpu_rdt\[18\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[15\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_123_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10825__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05965__A2 _02431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09998__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08903__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08116__B1 _03683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06390__A2 _02718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08945__S _04331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06142__A2 _02563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10205__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05576__S1 _01548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05420_ u_cpu.rf_ram.memory\[104\]\[3\] u_cpu.rf_ram.memory\[105\]\[3\] u_cpu.rf_ram.memory\[106\]\[3\]
+ u_cpu.rf_ram.memory\[107\]\[3\] _01615_ _01616_ _01909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_21_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08419__A1 _03788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05351_ u_cpu.rf_ram.memory\[88\]\[2\] u_cpu.rf_ram.memory\[89\]\[2\] u_cpu.rf_ram.memory\[90\]\[2\]
+ u_cpu.rf_ram.memory\[91\]\[2\] _01646_ _01603_ _01841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_119_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09092__A1 _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08070_ u_arbiter.i_wb_cpu_rdt\[13\] _03669_ _03678_ u_arbiter.i_wb_cpu_dbus_dat\[13\]
+ _03697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05282_ _01399_ _01772_ _01773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07642__A2 _03432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10355__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07021_ _02961_ _03081_ _03085_ _00418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09395__A2 _03798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05405__A1 _01601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08972_ _04346_ _01109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05956__A2 _01403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07923_ u_cpu.rf_ram.memory\[112\]\[3\] _03596_ _03600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09147__A2 _04439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06205__I0 _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07854_ _03547_ _03558_ _03562_ _00775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05708__A2 _02193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06905__A1 _02524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06805_ _02963_ _02955_ _02964_ _00323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07785_ u_cpu.rf_ram.memory\[34\]\[0\] _03520_ _03521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06381__A2 _02708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04997_ u_cpu.cpu.ctrl.o_ibus_adr\[20\] _01498_ _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09524_ _02475_ _02695_ _04663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08658__A1 u_arbiter.i_wb_cpu_ibus_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06736_ _02923_ _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06439__I _02501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08658__B2 u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09455_ u_cpu.rf_ram.memory\[24\]\[0\] _04625_ _04626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06667_ u_cpu.rf_ram.memory\[75\]\[1\] _02884_ _02886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06133__A2 _02551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05567__S1 _01580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08406_ _03816_ _03968_ _03975_ _03977_ _00912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_36_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05618_ _01609_ _02104_ _02105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09386_ u_cpu.cpu.decode.co_ebreak u_cpu.cpu.mem_bytecnt\[1\] u_cpu.cpu.mem_bytecnt\[0\]
+ _02337_ _04585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_24_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07881__A2 _02810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06598_ _02744_ _02844_ _02847_ _00233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05892__A1 _01370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08337_ u_cpu.cpu.immdec.imm24_20\[1\] _03798_ _03917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09083__A1 _02695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05549_ u_cpu.rf_ram.memory\[128\]\[4\] u_cpu.rf_ram.memory\[129\]\[4\] u_cpu.rf_ram.memory\[130\]\[4\]
+ u_cpu.rf_ram.memory\[131\]\[4\] _01687_ _01688_ _02037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__05319__S1 _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07633__A2 _03422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08268_ _03773_ _03858_ _03859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07219_ u_cpu.rf_ram.memory\[70\]\[1\] _03196_ _03198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08199_ _03797_ _03798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10848__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09386__A2 u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10230_ _00020_ io_in[4] u_cpu.rf_ram_if.rdata1\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07397__A1 _03157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10161_ _00607_ io_in[4] u_cpu.rf_ram.memory\[130\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10092_ _00538_ io_in[4] u_cpu.rf_ram.memory\[39\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05255__S0 _01590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06372__A2 _02708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10228__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08649__A1 _03551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10994_ _10994_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_43_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09310__A2 _04536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06124__A2 _02551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07321__A1 _03173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05558__S1 _01557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07872__A2 _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10378__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05883__A1 _01409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09074__A1 _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[69\] u_scanchain_local.module_data_in\[68\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[31\] u_scanchain_local.clk u_scanchain_local.module_data_in\[69\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_7_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09670__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07624__A2 _03422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08821__A1 _03825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06683__I0 _02573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10428_ _00861_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06812__I _02516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10359_ _00792_ io_in[4] u_cpu.rf_ram.memory\[8\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09129__A2 _04429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08188__I0 u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04920_ _01441_ _01442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08888__A1 _04284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05246__S0 _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05591__C _01628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04851_ u_cpu.cpu.decode.op21 _01371_ _01376_ _01377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_19_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07560__A1 _03357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06363__A2 _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07570_ _03349_ _03392_ _03395_ _00657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09301__A2 _04526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06521_ _02742_ _02801_ _02803_ _00200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06115__A2 _02541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05549__S1 _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09240_ _02584_ u_cpu.rf_ram.memory\[10\]\[2\] _04496_ _04499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06195__S _02603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06452_ _02573_ u_cpu.rf_ram.memory\[4\]\[0\] _02756_ _02757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07863__A2 _02821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05403_ _01597_ _01891_ _01892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09171_ u_cpu.rf_ram.memory\[108\]\[7\] _04449_ _04457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06383_ _02507_ _02708_ _02714_ _00151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09065__A1 _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08122_ _02539_ _02821_ _03730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05334_ u_cpu.rf_ram.memory\[100\]\[2\] u_cpu.rf_ram.memory\[101\]\[2\] u_cpu.rf_ram.memory\[102\]\[2\]
+ u_cpu.rf_ram.memory\[103\]\[2\] _01577_ _01549_ _01824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07615__A2 _03412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08812__A1 _03788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08812__B2 _03798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08053_ _03684_ _03685_ _00851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05265_ u_cpu.rf_ram.memory\[80\]\[1\] u_cpu.rf_ram.memory\[81\]\[1\] u_cpu.rf_ram.memory\[82\]\[1\]
+ u_cpu.rf_ram.memory\[83\]\[1\] _01545_ _01642_ _01756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_31_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07004_ u_cpu.rf_ram.memory\[54\]\[4\] _03071_ _03076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05721__S1 _01681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09368__A2 _04568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08415__I1 u_arbiter.i_wb_cpu_rdt\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05196_ _01668_ _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07379__A1 _03157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06051__A1 _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08955_ u_arbiter.i_wb_cpu_rdt\[22\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[6\]
+ _04331_ _04338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_102_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05782__B _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07906_ _03590_ _00799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08886_ _04280_ _04299_ _04300_ _01069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08879__A1 _04294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05237__S0 _01623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07837_ u_cpu.rf_ram.memory\[120\]\[5\] _03541_ _03552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09540__A2 _04664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06354__A2 _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07768_ _03343_ _03510_ _03511_ _00740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05073__I _01564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09507_ _04653_ _04654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06719_ u_cpu.rf_ram.memory\[67\]\[0\] _02914_ _02915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10520__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07699_ _03349_ _03465_ _03468_ _00713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06106__A2 _02541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07303__A1 _03173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09438_ _04468_ _04615_ _04616_ _01305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09693__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07854__A2 _03558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05865__A1 _01409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09056__A1 _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09369_ _01375_ _02306_ u_cpu.cpu.genblk3.csr.mcause3_0\[2\] _01385_ _04573_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_12_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10670__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07606__A2 _03412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08803__A1 _02312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08803__B2 _04010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05880__A4 _01375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08333__B _03913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04861__B _01386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05712__S1 _01652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09359__A2 _04556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06290__A1 _02517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05093__A2 _01584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10213_ _00659_ io_in[4] u_cpu.rf_ram.memory\[125\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10144_ _00590_ io_in[4] u_cpu.rf_ram.memory\[133\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07790__A1 _03349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06593__A2 _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10050__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10075_ _00521_ io_in[4] u_cpu.rf_ram.memory\[14\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05228__S0 _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09531__A2 _04664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07542__A1 _03357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06345__A2 _02686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05779__S1 _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06079__I _02527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_62_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10977_ _10977_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__09295__A1 _04474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07845__A2 _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05400__S0 _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09047__A1 _02682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[21\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05608__A1 _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08270__A2 _03802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05703__S1 _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05050_ _01541_ _01542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05084__A2 _01575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08022__A2 _02781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06033__A1 _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06584__A2 _02834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08740_ u_cpu.rf_ram.memory\[109\]\[4\] _04199_ _04204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05952_ u_cpu.rf_ram_if.rdata0\[2\] _01403_ _02425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05219__S0 _01578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09522__A2 _04654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04903_ _01403_ u_cpu.rf_ram_if.wtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_08671_ _04164_ _00990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__10543__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05883_ _01409_ _02363_ _02364_ _01372_ _02365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__05139__A3 _01588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06336__A2 _02686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07622_ _03347_ _03422_ _03424_ _00680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06918__S _03021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04898__A2 _01388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07553_ u_cpu.rf_ram.memory\[126\]\[3\] _03382_ _03386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08089__A2 _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06504_ u_cpu.rf_ram.memory\[16\]\[2\] _02791_ _02794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10693__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07484_ _02528_ _02893_ _03344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05847__A1 _01369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09223_ u_cpu.rf_ram.memory\[59\]\[2\] _04487_ _04490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06435_ _02744_ _02740_ _02745_ _00172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09038__A1 _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09154_ _04296_ _04439_ _04447_ _01190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06366_ _02512_ _02697_ _02704_ _00144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08105_ _03717_ _03718_ _03719_ _00869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05317_ _01601_ _01806_ _01605_ _01807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09085_ u_cpu.rf_ram.memory\[105\]\[0\] _04409_ _04410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05777__B _01564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06297_ _02487_ _02662_ _02664_ _00115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08261__A2 _03774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06272__A1 _02517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08036_ _03668_ _03669_ _03671_ _03672_ _00847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05248_ u_cpu.rf_ram.memory\[96\]\[1\] u_cpu.rf_ram.memory\[97\]\[1\] u_cpu.rf_ram.memory\[98\]\[1\]
+ u_cpu.rf_ram.memory\[99\]\[1\] _01602_ _01579_ _01739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_123_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09909__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09210__A1 _04480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10073__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05179_ u_cpu.rf_ram.memory\[68\]\[0\] u_cpu.rf_ram.memory\[69\]\[0\] u_cpu.rf_ram.memory\[70\]\[0\]
+ u_cpu.rf_ram.memory\[71\]\[0\] _01577_ _01549_ _01671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_104_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07072__I0 _02587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09987_ _00441_ io_in[4] u_cpu.rf_ram.memory\[15\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07772__A1 _03349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06575__A2 _02834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08938_ u_cpu.rf_ram.memory\[28\]\[6\] _04322_ _04329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09513__A2 _04654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08869_ u_cpu.rf_ram.memory\[94\]\[3\] _04282_ _04289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06327__A2 _02673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07524__A1 _03357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10900_ _01329_ io_in[4] u_cpu.rf_ram.memory\[98\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10831_ _01260_ io_in[4] u_cpu.rf_ram.memory\[111\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__04889__A2 _01414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09277__A1 _04474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04856__B _01381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10762_ _01191_ io_in[4] u_cpu.rf_ram.memory\[108\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[44\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09029__A1 _02810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10693_ _01122_ io_in[4] u_cpu.rf_ram.memory\[102\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10416__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05697__S0 _01623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09589__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08004__A2 _03636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09201__A1 _04474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07063__I0 _02599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10566__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06566__A2 _02823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10127_ _00573_ io_in[4] u_cpu.rf_ram.memory\[135\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09504__A2 _04644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10058_ _00504_ io_in[4] u_cpu.rf_ram.memory\[70\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06318__A2 _02673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07515__A1 u_cpu.rf_ram.memory\[128\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08712__B1 _04175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07818__A2 _03530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08953__S _04331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08491__A2 _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06220_ u_cpu.rf_ram.memory\[80\]\[3\] _02614_ _02618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05597__B _01416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06151_ u_cpu.rf_ram.memory\[20\]\[6\] _02563_ _02570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10096__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08243__A2 _03757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09440__A1 _04472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05102_ _01540_ _01594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06254__A1 u_cpu.cpu.immdec.imm11_7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05688__S0 _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06082_ u_cpu.rf_ram.memory\[21\]\[0\] _02530_ _02531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10909__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05033_ _01445_ _01527_ _01528_ u_arbiter.o_wb_cpu_adr\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09910_ _00364_ io_in[4] u_cpu.rf_ram.memory\[19\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06006__A1 _01386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09841_ _00295_ io_in[4] u_cpu.rf_ram.memory\[66\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06557__A2 _02823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07754__A1 _03349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08199__I _03797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09772_ _00226_ io_in[4] u_cpu.rf_ram.memory\[129\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06984_ u_cpu.rf_ram.memory\[55\]\[3\] _03061_ _03065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08723_ _04191_ _01386_ _04192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05935_ _02321_ u_cpu.rf_ram.rdata\[2\] _02414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06309__A2 _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08654_ _02305_ _02448_ _01428_ _04154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_39_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05866_ _01393_ _02348_ _02349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[67\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07605_ u_cpu.rf_ram.memory\[123\]\[2\] _03412_ _03415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09259__A1 _04474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08585_ _04114_ _00954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05797_ _02275_ _02277_ _02279_ _02281_ _01607_ _02282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_23_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07536_ _03351_ _03372_ _03376_ _00642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07809__A2 _03530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07467_ _02573_ u_cpu.rf_ram.memory\[12\]\[0\] _03334_ _03335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10439__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09206_ u_cpu.rf_ram.memory\[84\]\[4\] _04470_ _04479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07479__S _03334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06418_ _02502_ _02729_ _02734_ _00166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06493__A1 _01680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07398_ u_cpu.rf_ram.memory\[133\]\[1\] _03295_ _03297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09137_ _02475_ _02682_ _04438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09731__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06349_ _02517_ _02686_ _02694_ _00137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08234__A2 _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06245__A1 _02502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09068_ _04280_ _04399_ _04400_ _01151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10589__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06796__A2 _02955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08019_ _03648_ _03657_ _03658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11030_ _11030_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_89_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09881__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06548__A2 _02812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07745__A1 u_cpu.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05220__A2 _01710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08170__A1 _03765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05603__S0 _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06720__A2 _02914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10814_ _01243_ io_in[4] u_cpu.rf_ram.memory\[110\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10745_ _01174_ io_in[4] u_cpu.rf_ram.memory\[106\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08473__A2 _04016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06484__A1 _01408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10676_ _01105_ io_in[4] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[51\] u_scanchain_local.module_data_in\[50\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[13\] u_scanchain_local.clk u_scanchain_local.module_data_in\[51\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__08225__A2 _03778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09422__A1 _04472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07984__A1 _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06787__A2 _02944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.out_flop u_scanchain_local.module_data_in\[69\] u_scanchain_local.clk
+ u_scanchain_local.data_out_i vdd vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_110_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06539__A2 _02812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05720_ _02186_ _02205_ _01402_ _02206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_48_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09604__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08161__A1 _01435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05651_ _01562_ _02136_ _01565_ _02137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_64_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06711__A2 _02904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08370_ _03831_ _03773_ _03800_ _03940_ _03944_ _03945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_56_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05582_ _02062_ _02064_ _02066_ _02068_ _01607_ _02069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_143_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07321_ _03173_ _03245_ _03253_ _00550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_17_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09754__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06475__A1 u_arbiter.i_wb_cpu_dbus_dat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05278__A2 _01764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07252_ _02573_ u_cpu.rf_ram.memory\[14\]\[0\] _03215_ _03216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06203_ _02590_ u_cpu.rf_ram.memory\[7\]\[4\] _02603_ _02608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10731__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08216__A2 _03767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07183_ u_cpu.rf_ram.memory\[73\]\[1\] _03176_ _03178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06227__A1 _02512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06134_ _02517_ _02551_ _02559_ _00057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06778__A2 _02944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06065_ _02460_ u_cpu.cpu.o_wdata0 _02514_ _02515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10881__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05016_ u_arbiter.i_wb_cpu_dbus_adr\[24\] _01457_ _01516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07727__A1 _03359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09824_ _00278_ io_in[4] u_cpu.rf_ram.memory\[6\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05202__A2 _01693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10111__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09755_ _00209_ io_in[4] u_cpu.rf_ram.memory\[40\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06967_ _02961_ _03051_ _03055_ _00394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06950__A2 _03041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05918_ _02361_ _02396_ _02372_ _02399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_08706_ u_cpu.cpu.ctrl.o_ibus_adr\[23\] _04173_ _04175_ u_cpu.cpu.ctrl.o_ibus_adr\[24\]
+ _04183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09686_ _00140_ io_in[4] u_cpu.rf_ram.memory\[41\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06898_ _02963_ _03012_ _03017_ _00363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08637_ _04144_ _04145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05849_ _01370_ _02332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05505__A3 _01973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06702__A2 _02904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10261__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08593__S _04115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08568_ u_arbiter.i_wb_cpu_dbus_adr\[5\] u_arbiter.i_wb_cpu_dbus_adr\[4\] _02445_
+ _04106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05081__I _01548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07519_ u_cpu.rf_ram.memory\[128\]\[4\] _03362_ _03367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08499_ _03742_ _04027_ _03780_ _04060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08455__A2 _03797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10530_ _00963_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10461_ _00894_ io_in[4] u_cpu.cpu.decode.op22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08207__A2 _03798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09404__A1 _04472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07266__I0 _02599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10392_ _00825_ io_in[4] u_cpu.rf_ram.memory\[115\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07966__A1 _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06769__A2 _02934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11013_ _11013_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_133_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08766__I0 _02573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08768__S _04217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09627__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07194__A2 _03176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08391__A1 _03788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08391__B2 _03779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[30\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10604__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09777__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08694__A2 _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[45\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10754__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08446__A2 _02391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10728_ _01157_ io_in[4] u_cpu.rf_ram.memory\[79\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10659_ _01088_ io_in[4] u_cpu.rf_ram.memory\[28\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05432__A2 _01920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10134__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07709__A1 _03359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08757__I0 _02590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07870_ _03545_ _03568_ _03571_ _00782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08382__A1 _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07185__A2 _03176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06821_ u_cpu.rf_ram.memory\[63\]\[2\] _02972_ _02975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05815__S0 _01687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06932__A2 _03031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09540_ u_cpu.rf_ram.memory\[89\]\[7\] _04664_ _04672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10284__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06752_ _02754_ _02924_ _02932_ _00302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05703_ u_cpu.rf_ram.memory\[88\]\[6\] u_cpu.rf_ram.memory\[89\]\[6\] u_cpu.rf_ram.memory\[90\]\[6\]
+ u_cpu.rf_ram.memory\[91\]\[6\] _01646_ _01603_ _02189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_92_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09471_ _02577_ _02612_ _04634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06683_ _02573_ u_cpu.rf_ram.memory\[6\]\[0\] _02894_ _02895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_63_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08422_ u_cpu.cpu.immdec.imm30_25\[5\] _03954_ _03992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05634_ _01399_ _02120_ _02121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_58_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08353_ _03851_ _03926_ _03928_ _03929_ _03782_ _03930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_05565_ u_cpu.rf_ram.memory\[20\]\[5\] u_cpu.rf_ram.memory\[21\]\[5\] u_cpu.rf_ram.memory\[22\]\[5\]
+ u_cpu.rf_ram.memory\[23\]\[5\] _01572_ _01574_ _02052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08437__A2 _03988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07304_ _02695_ _02832_ _03244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08284_ _03756_ _03778_ _03779_ _03867_ _03851_ _03874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_05496_ _01609_ _01983_ _01984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06999__A2 _03071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07235_ u_cpu.rf_ram.memory\[143\]\[0\] _03206_ _03207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07166_ _03165_ _03159_ _03166_ _00482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07948__A1 _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06117_ _02469_ _02528_ _02550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08070__B1 _03678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07097_ _02967_ _03119_ _03126_ _00453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05423__A2 _01911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06620__A1 _02748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06048_ _02500_ _02501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10627__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05076__I _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08373__A1 _02305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09807_ _00261_ io_in[4] u_cpu.rf_ram.memory\[76\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05187__A1 _01657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07999_ u_cpu.rf_ram.memory\[33\]\[5\] _03636_ _03642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09738_ _00192_ io_in[4] u_cpu.rf_ram.memory\[16\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08125__A1 _03539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10777__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09669_ _00123_ io_in[4] u_cpu.rf_ram.memory\[44\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08676__A2 _04155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10007__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05679__C _01628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07100__A2 _02832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10513_ _00946_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10444_ _00877_ io_in[4] u_cpu.rf_ram.memory\[113\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10157__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08061__B1 _03678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10375_ _00808_ io_in[4] u_cpu.rf_ram.memory\[112\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05414__A2 _01902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[14\] u_arbiter.i_wb_cpu_rdt\[11\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[8\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_78_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08498__S _01437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05178__A1 _01667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06678__A1 _02752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05350__A1 _01398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08419__A2 _03786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05350_ _01398_ _01839_ _01840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08961__S _04331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09092__A2 _04409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05281_ u_cpu.rf_ram.memory\[136\]\[1\] u_cpu.rf_ram.memory\[137\]\[1\] u_cpu.rf_ram.memory\[138\]\[1\]
+ u_cpu.rf_ram.memory\[139\]\[1\] _01680_ _01681_ _01772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07020_ u_cpu.rf_ram.memory\[53\]\[3\] _03081_ _03085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06850__A1 _02969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08052__B1 _03678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05405__A2 _01893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06602__A1 _02748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08971_ u_arbiter.i_wb_cpu_rdt\[30\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[14\]
+ _04331_ _04346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09942__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07922_ _03545_ _03596_ _03599_ _00806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08355__A1 u_cpu.cpu.immdec.imm24_20\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07853_ u_cpu.rf_ram.memory\[118\]\[3\] _03558_ _03562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05169__A1 _01645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06905__A2 _02577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06804_ u_cpu.rf_ram.memory\[29\]\[4\] _02955_ _02964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07784_ _03519_ _03520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__04916__A1 _01437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04996_ _01443_ _01498_ _01499_ _01500_ u_arbiter.o_wb_cpu_adr\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_37_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09523_ _04484_ _04654_ _04662_ _01344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06735_ _02469_ _02626_ _02923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08658__A2 _04155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09454_ _04624_ _04625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_24_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06666_ _02738_ _02884_ _02885_ _00263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07330__A2 _03255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05617_ u_cpu.rf_ram.memory\[80\]\[5\] u_cpu.rf_ram.memory\[81\]\[5\] u_cpu.rf_ram.memory\[82\]\[5\]
+ u_cpu.rf_ram.memory\[83\]\[5\] _01590_ _01591_ _02104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08405_ u_cpu.cpu.immdec.imm30_25\[3\] _03949_ _03976_ u_cpu.cpu.immdec.imm30_25\[4\]
+ _03977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_52_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09385_ u_cpu.cpu.genblk3.csr.mie_mtie _04584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06597_ u_cpu.rf_ram.memory\[139\]\[2\] _02844_ _02847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07469__I0 _02581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08336_ _03915_ _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05548_ _01684_ _02035_ _01582_ _02036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09083__A2 _04197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08267_ _03831_ _03790_ _03858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05479_ u_cpu.rf_ram.memory\[16\]\[4\] u_cpu.rf_ram.memory\[17\]\[4\] u_cpu.rf_ram.memory\[18\]\[4\]
+ u_cpu.rf_ram.memory\[19\]\[4\] _01578_ _01580_ _01967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07218_ _03157_ _03196_ _03197_ _00503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08198_ _03796_ _03797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08969__I0 u_arbiter.i_wb_cpu_rdt\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08043__B1 _03678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07149_ _02596_ u_cpu.rf_ram.memory\[13\]\[6\] _03148_ _03155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09386__A3 u_cpu.cpu.mem_bytecnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07397__A2 _03295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10160_ _00606_ io_in[4] u_cpu.rf_ram.memory\[131\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10091_ _00537_ io_in[4] u_cpu.rf_ram.memory\[39\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08897__A2 _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05255__S1 _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10993_ _10993_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_90_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08649__A2 _04145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07321__A2 _03245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09815__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09074__A2 _04399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07085__A1 _02953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08821__A2 _03770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06832__A1 _02969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10427_ _00860_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09965__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07388__A2 _03285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10358_ _00791_ io_in[4] u_cpu.rf_ram.memory\[8\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05399__A1 _01589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10942__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10289_ _00722_ io_in[4] u_cpu.rf_ram.memory\[90\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08337__A1 u_cpu.cpu.immdec.imm24_20\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06199__I0 _02584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08888__A2 _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05246__S1 _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04850_ _01373_ _01375_ _01376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07560__A2 _03382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06520_ u_cpu.rf_ram.memory\[17\]\[1\] _02801_ _02803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07312__A2 _03245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10322__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06451_ _02561_ _02577_ _02756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05402_ u_cpu.rf_ram.memory\[60\]\[3\] u_cpu.rf_ram.memory\[61\]\[3\] u_cpu.rf_ram.memory\[62\]\[3\]
+ u_cpu.rf_ram.memory\[63\]\[3\] _01598_ _01573_ _01891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09170_ _04294_ _04449_ _04456_ _01197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06382_ u_cpu.rf_ram.memory\[43\]\[5\] _02708_ _02714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05874__A2 _02338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09065__A2 _02727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08121_ _03727_ _03678_ _03729_ _00875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05333_ _01594_ _01822_ _01416_ _01823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_30_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08812__A2 _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10472__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08052_ u_arbiter.i_wb_cpu_rdt\[7\] _03669_ _03678_ u_arbiter.i_wb_cpu_dbus_dat\[7\]
+ _03685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_31_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05264_ _01645_ _01754_ _01648_ _01755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05477__I2 u_cpu.rf_ram.memory\[22\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07003_ _02961_ _03071_ _03075_ _00410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05195_ _01571_ _01687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07379__A2 _03285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06051__A2 _02502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08954_ _04337_ _01100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08328__A1 _03773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07905_ _02587_ u_cpu.rf_ram.memory\[11\]\[3\] _03586_ _03590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08885_ u_cpu.rf_ram.memory\[95\]\[0\] _04299_ _04300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08879__A2 _04282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05237__S1 _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07836_ _02506_ _03551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07551__A2 _03382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07767_ u_cpu.rf_ram.memory\[35\]\[0\] _03510_ _03511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04979_ u_cpu.cpu.ctrl.o_ibus_adr\[13\] u_cpu.cpu.ctrl.o_ibus_adr\[12\] _01476_ _01487_
+ _01488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_25_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09506_ _02561_ _04197_ _04653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06718_ _02913_ _02914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07698_ u_cpu.rf_ram.memory\[91\]\[2\] _03465_ _03468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09838__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07303__A2 _03235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08500__A1 _03786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09437_ u_cpu.rf_ram.memory\[25\]\[0\] _04615_ _04616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06649_ u_cpu.rf_ram.memory\[76\]\[1\] _02874_ _02876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10815__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09368_ _02341_ _04568_ _04572_ _01279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09056__A2 _04389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09988__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08319_ _03779_ _03785_ _03900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09299_ _04478_ _04526_ _04531_ _01251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06814__A1 _02969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06290__A2 _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10212_ _00658_ io_in[4] u_cpu.rf_ram.memory\[125\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10143_ _00589_ io_in[4] u_cpu.rf_ram.memory\[133\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08319__A1 _03779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05250__B1 _01738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07790__A2 _03520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10074_ _00520_ io_in[4] u_cpu.rf_ram.memory\[14\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[7\] u_arbiter.i_wb_cpu_rdt\[4\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[1\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_47_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05228__S1 _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08776__S _04217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07542__A2 _03372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10345__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10976_ _10976_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__09295__A2 _04526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10495__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05856__A2 _01411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05400__S1 _01548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09047__A2 _04197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05608__A2 _02094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06805__A1 _02963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06281__A2 _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06033__A2 _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07230__A1 _03171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05883__B _01372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07781__A2 _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05951_ _01403_ _02322_ _02424_ _00008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05792__A1 _01645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04902_ _01399_ _01427_ _00025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_78_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08670_ u_cpu.cpu.ctrl.o_ibus_adr\[6\] _04155_ _04157_ u_cpu.cpu.ctrl.o_ibus_adr\[7\]
+ _04164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__05219__S1 _01580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05882_ _01369_ _01370_ _02364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_39_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07533__A2 _03372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08730__A1 _02660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07621_ u_cpu.rf_ram.memory\[38\]\[1\] _03422_ _03424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05544__A1 _02012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07552_ _03349_ _03382_ _03385_ _00649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10838__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09286__A2 _04516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06503_ _02742_ _02791_ _02793_ _00192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07297__A1 _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07483_ _02481_ _03343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05847__A2 _01390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06434_ u_cpu.rf_ram.memory\[50\]\[2\] _02740_ _02745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09222_ _04472_ _04487_ _04489_ _01216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09038__A2 _04379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09153_ u_cpu.rf_ram.memory\[83\]\[7\] _04439_ _04447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06365_ u_cpu.rf_ram.memory\[41\]\[6\] _02697_ _02704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08797__A1 _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08104_ u_arbiter.i_wb_cpu_rdt\[25\] _03653_ _03654_ u_arbiter.i_wb_cpu_dbus_dat\[25\]
+ _03719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05316_ u_cpu.rf_ram.memory\[56\]\[2\] u_cpu.rf_ram.memory\[57\]\[2\] u_cpu.rf_ram.memory\[58\]\[2\]
+ u_cpu.rf_ram.memory\[59\]\[2\] _01602_ _01579_ _01806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09084_ _04408_ _04409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05155__S0 _01646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06296_ u_cpu.rf_ram.memory\[45\]\[1\] _02662_ _02664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08035_ u_arbiter.i_wb_cpu_dbus_dat\[3\] _03664_ _03653_ _03672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05247_ _01636_ _01737_ _01738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06272__A2 _02641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10218__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08549__A1 _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05178_ _01667_ _01669_ _01670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09210__A2 _04470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09986_ _00440_ io_in[4] u_cpu.rf_ram.memory\[15\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07772__A2 _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10368__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08937_ _04292_ _04322_ _04328_ _01092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08868_ _02496_ _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09660__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07524__A2 _03362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07819_ _02481_ _03539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05535__A1 _01667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08799_ _03555_ _04227_ _04235_ _01047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10830_ _01259_ io_in[4] u_cpu.rf_ram.memory\[111\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09277__A2 _04516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10761_ _01190_ io_in[4] u_cpu.rf_ram.memory\[83\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05838__A2 _02321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09029__A2 _04197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10692_ _01121_ io_in[4] u_cpu.rf_ram.memory\[102\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08344__B _03797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06263__A2 _02641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05697__S1 _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[5\]_D u_arbiter.i_wb_cpu_rdt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09201__A2 _04470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07212__A1 _03171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07763__A2 _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10126_ _00572_ io_in[4] u_cpu.rf_ram.memory\[135\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10057_ _00503_ io_in[4] u_cpu.rf_ram.memory\[70\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07515__A2 _03362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05526__A1 _01398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09268__A2 _04506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07279__A1 _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10959_ _10959_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_17_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06150_ _02507_ _02563_ _02569_ _00063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_8_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09440__A2 _04615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05101_ _01589_ _01592_ _01593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07451__A1 _03157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06081_ _02529_ _02530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05688__S1 _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05032_ u_arbiter.i_wb_cpu_dbus_adr\[28\] _01457_ _01528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10510__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09840_ _00294_ io_in[4] u_cpu.rf_ram.memory\[67\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09683__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07754__A2 _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09771_ _00225_ io_in[4] u_cpu.rf_ram.memory\[129\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06983_ _02959_ _03061_ _03064_ _00401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08722_ _02343_ _01410_ _01378_ _04191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_100_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05934_ _02320_ _02412_ _02413_ _00015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_39_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10660__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05865_ _01409_ _02331_ _02334_ _02335_ _02347_ _02348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_08653_ _03555_ _04145_ _04153_ _00983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07604_ _03347_ _03412_ _03414_ _00672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_54_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05796_ _01614_ _02280_ _01654_ _02281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09259__A2 _04506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08584_ u_arbiter.i_wb_cpu_dbus_adr\[13\] u_arbiter.i_wb_cpu_dbus_adr\[12\] _02445_
+ _04114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_35_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07535_ u_cpu.rf_ram.memory\[127\]\[3\] _03372_ _03376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07466_ _02577_ _02671_ _03334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06417_ u_cpu.rf_ram.memory\[47\]\[4\] _02729_ _02734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09205_ _02501_ _04478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08219__B1 _03762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07690__A1 _01429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07397_ _03157_ _03295_ _03296_ _00583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10040__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09136_ _04296_ _04429_ _04437_ _01182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06348_ u_cpu.rf_ram.memory\[51\]\[7\] _02686_ _02694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09431__A2 _04605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06245__A2 _02628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09067_ u_cpu.rf_ram.memory\[79\]\[0\] _04399_ _04400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06279_ u_cpu.rf_ram.memory\[46\]\[2\] _02651_ _02654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05300__C _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05079__I _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07993__A2 _03636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08018_ u_arbiter.i_wb_cpu_dbus_dat\[0\] u_arbiter.i_wb_cpu_dbus_dat\[1\] _02774_
+ _03657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10190__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09195__A1 _04468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07745__A2 _03458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09969_ _00423_ io_in[4] u_cpu.rf_ram.memory\[52\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09498__A2 _04644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_u_scanchain_local.scan_flop\[11\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08170__A2 _03769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05603__S1 _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10813_ _01242_ io_in[4] u_cpu.rf_ram.memory\[110\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10744_ _01173_ io_in[4] u_cpu.rf_ram.memory\[106\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05698__B _01654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07681__A1 _01428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06484__A2 _01370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10675_ _01104_ io_in[4] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09422__A2 _04605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10533__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07433__A1 _03157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06236__A2 _02628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[44\] u_scanchain_local.module_data_in\[43\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[6\] u_scanchain_local.clk u_scanchain_local.module_data_in\[44\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_114_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07984__A2 _03626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05995__A1 u_cpu.cpu.bufreg.lsb\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09186__A1 _04292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10683__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08933__A1 _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10109_ _00555_ io_in[4] u_cpu.rf_ram.memory\[49\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11089_ _11089_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_110_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08161__A2 _03668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05650_ u_cpu.rf_ram.memory\[0\]\[6\] u_cpu.rf_ram.memory\[1\]\[6\] u_cpu.rf_ram.memory\[2\]\[6\]
+ u_cpu.rf_ram.memory\[3\]\[6\] _01556_ _01557_ _02136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_64_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05581_ _01601_ _02067_ _01605_ _02068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10063__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09110__A1 _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07320_ u_cpu.rf_ram.memory\[137\]\[7\] _03245_ _03253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05358__S0 _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07251_ _02577_ _02625_ _03215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06475__A2 _02770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07672__A1 _01428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10945__D u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06202_ _02607_ _00077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05401__B _01564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07182_ _03157_ _03176_ _03177_ _00487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09413__A2 _04595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06133_ u_cpu.rf_ram.memory\[18\]\[7\] _02551_ _02559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06227__A2 _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07975__A2 _03626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06064_ _02478_ u_cpu.rf_ram_if.wdata1_r\[7\] _02514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_133_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05015_ u_cpu.cpu.ctrl.o_ibus_adr\[24\] _01513_ _01515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_28_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07727__A2 _03475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[34\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08924__A1 _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09823_ _00277_ io_in[4] u_cpu.rf_ram.memory\[6\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09754_ _00208_ io_in[4] u_cpu.rf_ram.memory\[40\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06966_ u_cpu.rf_ram.memory\[56\]\[3\] _03051_ _03055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07842__I _02516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08705_ _04182_ _01006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_05917_ _02394_ _02397_ _02398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09685_ _00139_ io_in[4] u_cpu.rf_ram.memory\[41\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06897_ u_cpu.rf_ram.memory\[19\]\[4\] _03012_ _03017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08152__A2 _03751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10406__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08636_ _02528_ _02625_ _04144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_u_scanchain_local.scan_flop\[29\]_D u_arbiter.i_wb_cpu_rdt\[26\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_05848_ _01369_ _02309_ _02330_ _02331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09579__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08567_ _04105_ _00945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05910__A1 _01372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05779_ u_cpu.rf_ram.memory\[124\]\[7\] u_cpu.rf_ram.memory\[125\]\[7\] u_cpu.rf_ram.memory\[126\]\[7\]
+ u_cpu.rf_ram.memory\[127\]\[7\] _01545_ _01642_ _02264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09101__A1 _02638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07518_ _03351_ _03362_ _03366_ _00634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05349__S0 _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08498_ u_arbiter.i_wb_cpu_rdt\[18\] u_arbiter.i_wb_cpu_rdt\[2\] _01437_ _04059_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_11_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10556__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07449_ _03324_ _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_122_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10460_ _00893_ io_in[4] u_cpu.cpu.decode.op21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09404__A2 _04595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09119_ _02706_ _04197_ _04428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06218__A2 _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07415__A1 _03157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10391_ _00824_ io_in[4] u_cpu.rf_ram.memory\[115\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05426__B1 _01912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07966__A2 _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05521__S0 _01623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05977__A1 _02309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09168__A1 _04292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07718__A2 _03475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11012_ _11012_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_132_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08391__A2 _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05981__B _02445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10086__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06154__A1 _02517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10727_ _01156_ io_in[4] u_cpu.rf_ram.memory\[79\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10658_ _01087_ io_in[4] u_cpu.rf_ram.memory\[28\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05680__A3 _02165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10589_ _01019_ io_in[4] u_cpu.rf_ram.memory\[109\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07957__A2 _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[57\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05512__S0 _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05968__A1 u_cpu.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08959__S _04331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08906__A1 _04284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07709__A2 _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06820_ _02957_ _02972_ _02974_ _00328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10429__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05815__S1 _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06393__A1 _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06751_ u_cpu.rf_ram.memory\[66\]\[7\] _02924_ _02932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__04943__A2 _01457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09721__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08134__A2 _03731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09331__A1 _04474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05702_ _01398_ _02187_ _02188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06682_ _02577_ _02893_ _02894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09470_ _04484_ _04625_ _04633_ _01320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08421_ _03816_ _03985_ _03990_ _02768_ _03991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_24_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10579__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05633_ u_cpu.rf_ram.memory\[136\]\[5\] u_cpu.rf_ram.memory\[137\]\[5\] u_cpu.rf_ram.memory\[138\]\[5\]
+ u_cpu.rf_ram.memory\[139\]\[5\] _01680_ _01681_ _02120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_63_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05564_ _02044_ _02046_ _02048_ _02050_ _01568_ _02051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_08352_ _03890_ _03896_ _03851_ _03929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09871__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07303_ _03173_ _03235_ _03243_ _00542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08426__C _02438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05495_ u_cpu.rf_ram.memory\[40\]\[4\] u_cpu.rf_ram.memory\[41\]\[4\] u_cpu.rf_ram.memory\[42\]\[4\]
+ u_cpu.rf_ram.memory\[43\]\[4\] _01545_ _01642_ _01983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08283_ _03762_ _03828_ _03873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07234_ _03205_ _03206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09398__A1 _01428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07165_ u_cpu.rf_ram.memory\[72\]\[3\] _03159_ _03166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08442__B _03797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07948__A2 _03606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06116_ _02517_ _02541_ _02549_ _00049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08070__A1 u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07096_ u_cpu.rf_ram.memory\[142\]\[6\] _03119_ _03126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05959__A1 _01403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06047_ _02460_ u_cpu.rf_ram_if.wdata0_r\[4\] _02499_ _02500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06620__A2 _02854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05974__A4 _02438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08373__A2 _03947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09570__A1 _02769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09806_ _00260_ io_in[4] u_cpu.rf_ram.memory\[76\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_101_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07998_ _03549_ _03636_ _03641_ _00840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09737_ _00191_ io_in[4] u_cpu.rf_ram.memory\[16\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06949_ _02961_ _03041_ _03045_ _00386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04934__A2 _01443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08125__A2 _03731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09668_ _00122_ io_in[4] u_cpu.rf_ram.memory\[44\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08619_ u_arbiter.i_wb_cpu_dbus_adr\[30\] u_arbiter.i_wb_cpu_dbus_adr\[29\] _02372_
+ _04132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09599_ _00053_ io_in[4] u_cpu.rf_ram.memory\[18\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10512_ _00945_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10443_ _00876_ io_in[4] u_cpu.rf_ram.memory\[113\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08352__B _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07939__A2 _03606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08061__A1 u_arbiter.i_wb_cpu_rdt\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10374_ _00807_ io_in[4] u_cpu.rf_ram.memory\[112\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06611__A2 _02854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09744__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06375__A1 _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05178__A2 _01669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10721__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09313__A1 _04474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08116__A2 _03678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05216__B _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09894__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06678__A2 _02884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10871__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09202__I _02496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08246__C _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05280_ _01751_ _01770_ _01402_ _01771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10101__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06850__A2 _02982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08052__A1 u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06602__A2 _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08970_ _04345_ _01108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10251__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07921_ u_cpu.rf_ram.memory\[112\]\[2\] _03596_ _03599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08355__A2 _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07852_ _03545_ _03558_ _03561_ _00774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06366__A1 _02512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05169__A2 _01660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06803_ _02501_ _02963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07783_ _02469_ _02639_ _03519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04995_ u_arbiter.i_wb_cpu_dbus_adr\[19\] _01442_ _01500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08107__A2 _03678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09522_ u_cpu.rf_ram.memory\[100\]\[7\] _04654_ _04662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05126__B _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06734_ _02754_ _02914_ _02922_ _00294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05841__S _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07866__A1 _03539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09453_ _02528_ _02810_ _04624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06669__A2 _02884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06665_ u_cpu.rf_ram.memory\[75\]\[0\] _02884_ _02885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08404_ _02305_ _03796_ _03947_ _03976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05616_ _01645_ _02102_ _01648_ _02103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09384_ _04583_ _01284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06596_ _02742_ _02844_ _02846_ _00232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08335_ _03796_ _03914_ _03915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_71_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08815__B1 _03809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05547_ u_cpu.rf_ram.memory\[140\]\[4\] u_cpu.rf_ram.memory\[141\]\[4\] u_cpu.rf_ram.memory\[142\]\[4\]
+ u_cpu.rf_ram.memory\[143\]\[4\] _01680_ _01681_ _02035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_137_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09617__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08266_ _03761_ _03828_ _03857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07094__A2 _03119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05478_ _01570_ _01965_ _01966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07217_ u_cpu.rf_ram.memory\[70\]\[0\] _03196_ _03197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05796__B _01654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06841__A2 _02982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08197_ u_arbiter.i_wb_cpu_ack _01431_ _03795_ _03796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_106_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04852__A1 _01372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06471__I _02767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08043__A1 u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07148_ _03154_ _00476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09386__A4 _02337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09767__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07079_ _03116_ _00445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08599__S _04115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05087__I _01547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[44\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10090_ _00536_ io_in[4] u_cpu.rf_ram.memory\[39\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10744__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[59\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10992_ _10992_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__10894__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10124__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08282__A1 _03762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07085__A2 _03119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06832__A2 _02972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10274__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10426_ _00859_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10357_ _00790_ io_in[4] u_cpu.rf_ram.memory\[8\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06596__A1 _02742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10288_ _00721_ io_in[4] u_cpu.rf_ram.memory\[90\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08337__A2 _03798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06899__A2 _03012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05020__A1 u_arbiter.i_wb_cpu_dbus_adr\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07848__A1 _03539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08257__B _03831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06450_ _02754_ _02740_ _02755_ _00177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05401_ _01594_ _01889_ _01564_ _01890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06381_ _02502_ _02708_ _02713_ _00150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05332_ u_cpu.rf_ram.memory\[104\]\[2\] u_cpu.rf_ram.memory\[105\]\[2\] u_cpu.rf_ram.memory\[106\]\[2\]
+ u_cpu.rf_ram.memory\[107\]\[2\] _01615_ _01616_ _01822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10617__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08120_ u_arbiter.i_wb_cpu_rdt\[31\] _02781_ _03718_ _02325_ _03729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_119_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08273__A1 _03800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08273__B2 _03761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05263_ u_cpu.rf_ram.memory\[88\]\[1\] u_cpu.rf_ram.memory\[89\]\[1\] u_cpu.rf_ram.memory\[90\]\[1\]
+ u_cpu.rf_ram.memory\[91\]\[1\] _01646_ _01603_ _01754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08051_ u_arbiter.i_wb_cpu_dbus_dat\[8\] _03683_ _03684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06823__A2 _02972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07002_ u_cpu.rf_ram.memory\[54\]\[3\] _03071_ _03075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08025__A1 u_arbiter.i_wb_cpu_dbus_dat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05194_ _01684_ _01685_ _01582_ _01686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10767__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08953_ u_arbiter.i_wb_cpu_rdt\[21\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[5\]
+ _04331_ _04337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07904_ _03589_ _00798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08884_ _04298_ _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_111_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06339__A1 _02492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07835_ _03549_ _03541_ _03550_ _00768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07000__A2 _03071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07766_ _03509_ _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07139__I0 _02581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04978_ u_cpu.cpu.ctrl.o_ibus_adr\[15\] u_cpu.cpu.ctrl.o_ibus_adr\[14\] _01487_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_72_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10147__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09505_ _04484_ _04644_ _04652_ _01336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06717_ _02626_ _02682_ _02913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07697_ _03347_ _03465_ _03467_ _00712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08500__A2 _03860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09436_ _04614_ _04615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06648_ _02738_ _02874_ _02875_ _00255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06511__A1 _02750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09367_ _04568_ _04571_ _04572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06579_ u_cpu.rf_ram.memory\[129\]\[2\] _02834_ _02837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10297__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08318_ _03898_ _03899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_123_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08264__A1 _01381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09298_ u_cpu.rf_ram.memory\[86\]\[4\] _04526_ _04531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08249_ _03841_ _03842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06814__A2 _02955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10211_ _00657_ io_in[4] u_cpu.rf_ram.memory\[125\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06578__A1 _02742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10142_ _00588_ io_in[4] u_cpu.rf_ram.memory\[133\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08319__A2 _03785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10073_ _00519_ io_in[4] u_cpu.rf_ram.memory\[14\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06750__A1 _02752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10975_ _10975_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_44_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09932__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08255__A1 _03752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08255__B2 _03763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05069__A1 _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06805__A2 _02955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08007__A1 _02305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08558__A2 _04094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10409_ _00842_ io_in[4] u_cpu.rf_ram.memory\[33\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06569__A1 _02752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07230__A2 _03196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05241__A1 _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05092__I1 u_cpu.rf_ram.memory\[29\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05950_ u_cpu.rf_ram_if.rdata0\[1\] _01403_ _02424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08967__S _04331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04901_ _01406_ _01418_ _01422_ _01426_ _01427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_66_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05881_ u_cpu.cpu.branch_op _02313_ _02363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_38_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08730__A2 _04197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07620_ _03343_ _03422_ _03423_ _00679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07551_ u_cpu.rf_ram.memory\[126\]\[2\] _03382_ _03385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06502_ u_cpu.rf_ram.memory\[16\]\[1\] _02791_ _02793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07297__A2 _03235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08494__A1 _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07482_ _03342_ _00622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09221_ u_cpu.rf_ram.memory\[59\]\[1\] _04487_ _04489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06433_ _02491_ _02744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09152_ _04294_ _04439_ _04446_ _01189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06364_ _02507_ _02697_ _02703_ _00143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08103_ _02781_ _03648_ _03718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08797__A2 _04227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05315_ _01597_ _01804_ _01805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06295_ _02482_ _02662_ _02663_ _00114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09083_ _02695_ _04197_ _04408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05155__S1 _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08034_ u_arbiter.i_wb_cpu_dbus_dat\[4\] _02774_ _03648_ _03670_ _03671_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05246_ u_cpu.rf_ram.memory\[100\]\[1\] u_cpu.rf_ram.memory\[101\]\[1\] u_cpu.rf_ram.memory\[102\]\[1\]
+ u_cpu.rf_ram.memory\[103\]\[1\] _01598_ _01573_ _01737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_128_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05480__A1 _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08549__A2 _04094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05177_ u_cpu.rf_ram.memory\[64\]\[0\] u_cpu.rf_ram.memory\[65\]\[0\] u_cpu.rf_ram.memory\[66\]\[0\]
+ u_cpu.rf_ram.memory\[67\]\[0\] _01571_ _01668_ _01669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_143_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07221__A2 _03196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09985_ _00439_ io_in[4] u_cpu.rf_ram.memory\[15\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05232__A1 _01609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08936_ u_cpu.rf_ram.memory\[28\]\[5\] _04322_ _04328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09805__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08867_ _04286_ _04282_ _04287_ _01063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07818_ _03359_ _03530_ _03538_ _00763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08798_ u_cpu.rf_ram.memory\[93\]\[7\] _04227_ _04235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06732__A1 _02752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05535__A2 _02022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07749_ u_cpu.rf_ram.memory\[92\]\[0\] _03500_ _03501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09955__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10760_ _01189_ io_in[4] u_cpu.rf_ram.memory\[83\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07288__A2 _03235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05299__A1 _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09419_ u_cpu.rf_ram.memory\[26\]\[0\] _04605_ _04606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10691_ _01120_ io_in[4] u_cpu.rf_ram.memory\[102\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10932__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08237__A1 _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08788__A2 _04227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06799__A1 _02959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07460__A2 _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05471__A1 _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07212__A2 _03186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10312__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05223__A1 _01589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10125_ _00571_ io_in[4] u_cpu.rf_ram.memory\[135\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06971__A1 _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10056_ _00502_ io_in[4] u_cpu.rf_ram.memory\[71\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_u_scanchain_local.scan_flop\[8\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08712__A2 _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10462__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08586__I _02372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05526__A2 _02013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08476__A1 _03788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07279__A2 _03225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10958_ _10958_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_32_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10889_ _01318_ io_in[4] u_cpu.rf_ram.memory\[24\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08228__A1 _01374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05100_ u_cpu.rf_ram.memory\[52\]\[0\] u_cpu.rf_ram.memory\[53\]\[0\] u_cpu.rf_ram.memory\[54\]\[0\]
+ u_cpu.rf_ram.memory\[55\]\[0\] _01590_ _01591_ _01592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_06080_ _02524_ _02528_ _02529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07451__A2 _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05031_ u_cpu.cpu.ctrl.o_ibus_adr\[28\] _01526_ _01527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__05462__A1 _01399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09828__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08400__A1 _01436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07203__A2 _03186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05214__A1 _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09770_ _00224_ io_in[4] u_cpu.rf_ram.memory\[129\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06982_ u_cpu.rf_ram.memory\[55\]\[2\] _03061_ _03064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10805__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08721_ _04190_ _01014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05933_ _02320_ u_cpu.rf_ram_if.rdata1\[1\] _02413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09978__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08652_ u_cpu.rf_ram.memory\[30\]\[7\] _04145_ _04153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05864_ _02336_ _02324_ _02340_ u_cpu.cpu.genblk3.csr.mstatus_mie _02346_ _02347_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_66_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06714__A1 _02752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07603_ u_cpu.rf_ram.memory\[123\]\[1\] _03412_ _03414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08583_ _04113_ _00953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05795_ u_cpu.rf_ram.memory\[84\]\[7\] u_cpu.rf_ram.memory\[85\]\[7\] u_cpu.rf_ram.memory\[86\]\[7\]
+ u_cpu.rf_ram.memory\[87\]\[7\] _01555_ _01652_ _02280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10955__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07534_ _03349_ _03372_ _03375_ _00641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08467__A1 _03890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07465_ _03173_ _03325_ _03333_ _00614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09204_ _04476_ _04470_ _04477_ _01210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06416_ _02497_ _02729_ _02733_ _00165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08219__A1 _01372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08219__B2 _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07396_ u_cpu.rf_ram.memory\[133\]\[0\] _03295_ _03296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09135_ u_cpu.rf_ram.memory\[107\]\[7\] _04429_ _04437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06347_ _02512_ _02686_ _02693_ _00136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09066_ _04398_ _04399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06278_ _02487_ _02651_ _02653_ _00107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07442__A2 _03315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10335__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05453__A1 _01636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08017_ u_arbiter.i_wb_cpu_dbus_dat\[2\] _02774_ _03656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05229_ _01601_ _01719_ _01605_ _01720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09195__A2 _04470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05205__A1 _01542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10485__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09968_ _00422_ io_in[4] u_cpu.rf_ram.memory\[53\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06953__A1 _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08919_ u_cpu.cpu.bufreg.i_sh_signed _03798_ _04318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09899_ _00353_ io_in[4] u_cpu.rf_ram.memory\[60\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05823__I _01409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08339__C _03855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10812_ _01241_ io_in[4] u_cpu.rf_ram.memory\[110\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10743_ _01172_ io_in[4] u_cpu.rf_ram.memory\[106\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06484__A3 _02779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10674_ _01103_ io_in[4] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05692__A1 _01589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08630__A1 u_cpu.cpu.bufreg.lsb\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08091__C1 _03676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07433__A2 _03315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05444__A1 _01553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_scanchain_local.scan_flop\[37\] u_scanchain_local.module_data_in\[36\] io_in[3]
+ u_arbiter.i_wb_cpu_dbus_dat\[31\] u_scanchain_local.clk u_scanchain_local.module_data_in\[37\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__05995__A2 u_cpu.cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10828__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09186__A2 _04459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07197__A1 _02602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08933__A2 _04322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10108_ _00554_ io_in[4] u_cpu.rf_ram.memory\[49\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11088_ _11088_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10039_ _00485_ io_in[4] u_cpu.rf_ram.memory\[72\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09205__I _02501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10208__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05580_ u_cpu.rf_ram.memory\[56\]\[5\] u_cpu.rf_ram.memory\[57\]\[5\] u_cpu.rf_ram.memory\[58\]\[5\]
+ u_cpu.rf_ram.memory\[59\]\[5\] _01602_ _01579_ _02067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_32_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09110__A2 _04419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07121__A1 _02953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05358__S1 _01668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07250_ _03173_ _03206_ _03214_ _00518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10358__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05683__A1 _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06201_ _02587_ u_cpu.rf_ram.memory\[7\]\[3\] _02603_ _02607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07181_ u_cpu.rf_ram.memory\[73\]\[0\] _03176_ _03177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09650__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06132_ _02512_ _02551_ _02558_ _00056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07424__A2 _03305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06063_ _02477_ _02512_ _02513_ _00032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05014_ _01443_ _01511_ _01513_ _01514_ u_arbiter.o_wb_cpu_adr\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__09177__A2 _04459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07188__A1 _03165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09822_ _00276_ io_in[4] u_cpu.rf_ram.memory\[6\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08924__A2 _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06935__A1 _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05294__S0 _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09753_ _00207_ io_in[4] u_cpu.rf_ram.memory\[40\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06965_ _02959_ _03051_ _03054_ _00393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08704_ u_cpu.cpu.ctrl.o_ibus_adr\[22\] _04173_ _04175_ u_cpu.cpu.ctrl.o_ibus_adr\[23\]
+ _04182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05916_ u_cpu.cpu.mem_bytecnt\[1\] _02395_ _02396_ _02397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09684_ _00138_ io_in[4] u_cpu.rf_ram.memory\[41\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06896_ _02961_ _03012_ _03016_ _00362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08635_ _02431_ _04139_ _04143_ _00975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05847_ _01369_ _01390_ _02330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08566_ u_arbiter.i_wb_cpu_dbus_adr\[4\] u_arbiter.i_wb_cpu_dbus_adr\[3\] _02445_
+ _04105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_14_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05778_ _02256_ _02258_ _02260_ _02262_ _01628_ _02263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_70_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05910__A2 _02313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09101__A2 _04197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07517_ u_cpu.rf_ram.memory\[128\]\[3\] _03362_ _03366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08497_ _04016_ _04056_ _04057_ _04058_ _00922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_74_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05349__S1 _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07448_ _02469_ _02832_ _03324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07663__A2 _03442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05674__A1 _01397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07379_ _03157_ _03285_ _03286_ _00575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09118_ _04296_ _04419_ _04427_ _01174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10390_ _00823_ io_in[4] u_cpu.rf_ram.memory\[115\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07415__A2 _03305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09049_ u_cpu.rf_ram.memory\[99\]\[0\] _04389_ _04390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05521__S1 _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09168__A2 _04449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07179__A1 _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11011_ _11011_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__08915__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05285__S0 _01687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04878__B _01403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09340__A2 _04546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07351__A1 _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06154__A2 _02563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10500__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07103__A1 _02953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09673__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05502__B _01626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10726_ _01155_ io_in[4] u_cpu.rf_ram.memory\[79\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05665__A1 _01540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10657_ _01086_ io_in[4] u_cpu.cpu.genblk1.align.ctrl_misal vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05221__C _01426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10650__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07406__A2 _03295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10588_ _01018_ io_in[4] u_cpu.rf_ram.memory\[109\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05417__A1 _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05512__S1 _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05968__A2 _02433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09159__A2 _04449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08906__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05276__S0 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08119__B1 _03683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07590__A1 _03351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06393__A2 _02718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10030__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06750_ _02752_ _02924_ _02931_ _00301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05701_ u_cpu.rf_ram.memory\[92\]\[6\] u_cpu.rf_ram.memory\[93\]\[6\] u_cpu.rf_ram.memory\[94\]\[6\]
+ u_cpu.rf_ram.memory\[95\]\[6\] _01610_ _01611_ _02187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09331__A2 _04546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06681_ _02468_ _02523_ _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_63_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06145__A2 _02563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08390__I0 u_arbiter.i_wb_cpu_rdt\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08420_ _03987_ _03989_ _03906_ _03990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_64_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05632_ _02099_ _02118_ _01402_ _02119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10180__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08351_ _03776_ _03923_ _03927_ _03826_ _03928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05563_ _01562_ _02049_ _01565_ _02050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08142__I0 u_arbiter.i_wb_cpu_rdt\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07302_ u_cpu.rf_ram.memory\[39\]\[7\] _03235_ _03243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08282_ _03762_ _03868_ _03871_ _03872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08842__A1 _03539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07645__A2 _03432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05494_ _01975_ _01977_ _01979_ _01981_ _01607_ _01982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__05656__A1 _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07233_ _02727_ _02832_ _03205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07164_ _02496_ _03165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05408__A1 _01609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06115_ u_cpu.rf_ram.memory\[81\]\[7\] _02541_ _02549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06456__I0 _02584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08070__A2 _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07095_ _02965_ _03119_ _03125_ _00452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06046_ _02478_ u_cpu.rf_ram_if.wdata1_r\[4\] _02499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_99_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05267__S0 _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09805_ _00259_ io_in[4] u_cpu.rf_ram.memory\[76\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07997_ u_cpu.rf_ram.memory\[33\]\[4\] _03636_ _03641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07581__A1 _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06384__A2 _02708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09736_ _00190_ io_in[4] u_cpu.raddr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06948_ u_cpu.rf_ram.memory\[57\]\[3\] _03041_ _03045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09322__A2 _04536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09667_ _00121_ io_in[4] u_cpu.rf_ram.memory\[45\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10523__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06879_ u_cpu.rf_ram.memory\[60\]\[4\] _03002_ _03007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07333__A1 _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08618_ _04131_ _00970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09696__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09598_ _00052_ io_in[4] u_cpu.rf_ram.memory\[18\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08549_ _03543_ _04094_ _04096_ _00936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09086__A1 _04280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05322__B _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10673__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08833__A1 _03773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05647__A1 _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10511_ _00944_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06695__I0 _02596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10442_ _00875_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10373_ _00806_ io_in[4] u_cpu.rf_ram.memory\[112\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08061__A2 _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09010__A1 _04296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10053__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09561__A2 _04683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07572__A1 _03351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06375__A2 _02708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09313__A2 _04536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06127__A2 _02551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07875__A2 _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05886__A1 u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07627__A2 _03422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[24\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08824__A1 u_cpu.cpu.immdec.imm11_7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08824__B2 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05638__A1 _01399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10709_ _01138_ io_in[4] u_cpu.rf_ram.memory\[104\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08052__A2 _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06063__A1 _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05497__S0 _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07920_ _03543_ _03596_ _03598_ _00805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05810__A1 _01399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07851_ u_cpu.rf_ram.memory\[118\]\[2\] _03558_ _03561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09552__A2 _04674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10546__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07563__A1 _02660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06366__A2 _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06802_ _02961_ _02955_ _02962_ _00322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07782_ _03359_ _03510_ _03518_ _00747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_7_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04994_ u_cpu.cpu.ctrl.o_ibus_adr\[19\] _01495_ _01499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09521_ _04482_ _04654_ _04661_ _01343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09304__A2 _04526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06733_ u_cpu.rf_ram.memory\[67\]\[7\] _02914_ _02922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07315__A1 _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09452_ _04484_ _04615_ _04623_ _01312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10696__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06664_ _02883_ _02884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07866__A2 _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08403_ _03812_ _03971_ _03974_ _03975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_51_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05615_ u_cpu.rf_ram.memory\[88\]\[5\] u_cpu.rf_ram.memory\[89\]\[5\] u_cpu.rf_ram.memory\[90\]\[5\]
+ u_cpu.rf_ram.memory\[91\]\[5\] _01646_ _01603_ _02102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08437__C _03801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09383_ u_cpu.cpu.genblk3.csr.mstatus_mie u_cpu.cpu.genblk3.csr.mstatus_mpie _04565_
+ _04583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09068__A1 _04280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06595_ u_cpu.rf_ram.memory\[139\]\[1\] _02844_ _02846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08334_ _02436_ _02313_ _01376_ _02305_ _03914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_05546_ _01399_ _02033_ _02034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08815__A1 _03973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08815__B2 _03757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05629__A1 _01553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08265_ u_arbiter.i_wb_cpu_rdt\[21\] u_arbiter.i_wb_cpu_rdt\[5\] _01437_ _03856_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08291__A2 _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05477_ u_cpu.rf_ram.memory\[20\]\[4\] u_cpu.rf_ram.memory\[21\]\[4\] u_cpu.rf_ram.memory\[22\]\[4\]
+ u_cpu.rf_ram.memory\[23\]\[4\] _01572_ _01574_ _01965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_137_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07216_ _03195_ _03196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08196_ _02765_ u_arbiter.i_wb_cpu_ibus_adr\[1\] _03795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04852__A2 _01374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07147_ _02593_ u_cpu.rf_ram.memory\[13\]\[5\] _03148_ _03154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10076__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08043__A2 _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05488__S0 _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07078_ _02596_ u_cpu.rf_ram.memory\[15\]\[6\] _03109_ _03116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_126_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05801__A1 _01553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06029_ _02460_ u_cpu.rf_ram_if.wdata0_r\[1\] _02484_ _02485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_133_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07554__A1 _03351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06357__A2 _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05317__B _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09719_ _00173_ io_in[4] u_cpu.rf_ram.memory\[50\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10991_ _10991_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__06109__A2 _02541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08628__B _02338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07857__A2 _03558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[47\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07609__A2 _03412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10419__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10425_ _00858_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09711__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08034__A2 _02774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06045__A1 _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05479__S0 _01578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10356_ _00789_ io_in[4] u_cpu.rf_ram.memory\[8\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10569__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[54\]_SI u_arbiter.o_wb_cpu_adr\[16\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06596__A2 _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10287_ _00720_ io_in[4] u_cpu.rf_ram.memory\[90\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09861__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09534__A2 _04664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07545__A1 _02625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06348__A2 _02686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05020__A2 _01457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07848__A2 _03558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05859__A1 _02311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06520__A2 _02801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05400_ u_cpu.rf_ram.memory\[48\]\[3\] u_cpu.rf_ram.memory\[49\]\[3\] u_cpu.rf_ram.memory\[50\]\[3\]
+ u_cpu.rf_ram.memory\[51\]\[3\] _01544_ _01548_ _01889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_06380_ u_cpu.rf_ram.memory\[43\]\[4\] _02708_ _02713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05331_ _01597_ _01820_ _01821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10099__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09470__A1 _04484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06284__A1 _02502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08050_ _03676_ _03683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05262_ _01398_ _01752_ _01753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07001_ _02959_ _03071_ _03074_ _00409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08025__A2 u_arbiter.i_wb_cpu_dbus_dat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05193_ u_cpu.rf_ram.memory\[140\]\[0\] u_cpu.rf_ram.memory\[141\]\[0\] u_cpu.rf_ram.memory\[142\]\[0\]
+ u_cpu.rf_ram.memory\[143\]\[0\] _01680_ _01681_ _01685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09222__A1 _04472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05188__I _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06587__A2 _02834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08952_ _04336_ _01099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07903_ _02584_ u_cpu.rf_ram.memory\[11\]\[2\] _03586_ _03589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08883_ _02475_ _02727_ _04298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07536__A1 _03351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06339__A2 _02686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07834_ u_cpu.rf_ram.memory\[120\]\[4\] _03541_ _03550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07765_ _02639_ _02682_ _03509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04977_ u_cpu.cpu.ctrl.o_ibus_adr\[14\] _01481_ u_cpu.cpu.ctrl.o_ibus_adr\[15\] _01486_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_72_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09504_ u_cpu.rf_ram.memory\[98\]\[7\] _04644_ _04652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06716_ _02754_ _02904_ _02912_ _00286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07696_ u_cpu.rf_ram.memory\[91\]\[1\] _03465_ _03467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09435_ _02528_ _02695_ _04614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06647_ u_cpu.rf_ram.memory\[76\]\[0\] _02874_ _02875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06511__A2 _02791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09366_ _04569_ _04570_ _04571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06683__S _02894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06578_ _02742_ _02834_ _02836_ _00224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_127_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08317_ _03831_ _03776_ _03898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05529_ u_cpu.rf_ram.memory\[80\]\[4\] u_cpu.rf_ram.memory\[81\]\[4\] u_cpu.rf_ram.memory\[82\]\[4\]
+ u_cpu.rf_ram.memory\[83\]\[4\] _01590_ _01591_ _02017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09297_ _04476_ _04526_ _04530_ _01250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08264__A2 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09734__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08248_ _03757_ _03759_ _03819_ _03841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_119_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10711__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09213__A1 _04482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08179_ _03776_ _03778_ _03779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05098__I _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10210_ _00656_ io_in[4] u_cpu.rf_ram.memory\[125\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06027__A1 _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09884__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08811__I1 u_cpu.cpu.immdec.imm11_7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06578__A2 _02834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10141_ _00587_ io_in[4] u_cpu.rf_ram.memory\[133\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10861__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09516__A2 _04654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10072_ _00518_ io_in[4] u_cpu.rf_ram.memory\[143\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07527__A1 _02727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05002__A2 _01457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05633__S0 _01680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06750__A2 _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10974_ _10974_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_62_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06502__A2 _02791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10241__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08255__A2 _03770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[67\] u_scanchain_local.module_data_in\[66\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[29\] u_scanchain_local.clk u_scanchain_local.module_data_in\[67\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__09452__A1 _04484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07488__I _02486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06266__A1 _02502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05069__A2 _01560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04905__I _01428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10391__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09204__A1 _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10408_ _00841_ io_in[4] u_cpu.rf_ram.memory\[33\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07066__I0 _02573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06569__A2 _02823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10339_ _00772_ io_in[4] u_cpu.rf_ram.memory\[118\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09208__I _02506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05241__A2 _01703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07518__A1 _03351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08566__I0 u_arbiter.i_wb_cpu_dbus_adr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04900_ _01425_ _01426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_78_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05880_ _01384_ u_cpu.cpu.state.init_done _01385_ _01375_ _02362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_61_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09607__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08191__A1 _03754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05624__S0 _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06741__A2 _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07550_ _03347_ _03382_ _03384_ _00648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_93_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06501_ _02738_ _02791_ _02792_ _00191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07481_ _02599_ u_cpu.rf_ram.memory\[12\]\[7\] _03334_ _03342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_59_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09757__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09220_ _04468_ _04487_ _04488_ _01215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06432_ _02742_ _02740_ _02743_ _00171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[43\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09151_ u_cpu.rf_ram.memory\[83\]\[6\] _04439_ _04446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10734__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06363_ u_cpu.rf_ram.memory\[41\]\[5\] _02697_ _02703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08246__A2 _03802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08102_ u_arbiter.i_wb_cpu_dbus_dat\[26\] _03717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05314_ u_cpu.rf_ram.memory\[60\]\[2\] u_cpu.rf_ram.memory\[61\]\[2\] u_cpu.rf_ram.memory\[62\]\[2\]
+ u_cpu.rf_ram.memory\[63\]\[2\] _01598_ _01573_ _01804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_120_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09082_ _04296_ _04399_ _04407_ _01158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06294_ u_cpu.rf_ram.memory\[45\]\[0\] _02662_ _02663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08033_ _02774_ _02775_ _03670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05245_ _01594_ _01735_ _01416_ _01736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_u_scanchain_local.scan_flop\[58\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06009__A1 _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07057__I0 _02590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10884__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05176_ _01548_ _01668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09984_ _00438_ io_in[4] u_cpu.rf_ram.memory\[9\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05232__A2 _01722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05083__I2 u_cpu.rf_ram.memory\[22\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10114__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08935_ _04290_ _04322_ _04327_ _01091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07509__A1 _02612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08706__B1 _04175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06980__A2 _03061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08866_ u_cpu.rf_ram.memory\[94\]\[2\] _04282_ _04287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08182__A1 _03774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05615__S0 _01646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07817_ u_cpu.rf_ram.memory\[117\]\[7\] _03530_ _03538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08797_ _03553_ _04227_ _04234_ _01046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08309__I0 u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06732__A2 _02914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10264__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07748_ _03499_ _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_77_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07679_ u_cpu.cpu.mem_bytecnt\[0\] _03454_ _03456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08485__A2 _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06496__A1 _01681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09418_ _04604_ _04605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10690_ _01119_ io_in[4] u_cpu.rf_ram.memory\[102\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09349_ _04474_ _04556_ _04559_ _01273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09434__A1 _04484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07996__A1 _03547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06799__A2 _02955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05471__A2 _01958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06420__A1 _02507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10124_ _00570_ io_in[4] u_cpu.rf_ram.memory\[135\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05223__A2 _01713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06971__A2 _03051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10055_ _00501_ io_in[4] u_cpu.rf_ram.memory\[71\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10607__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07920__A1 _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06723__A2 _02914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10757__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10957_ _10957_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_90_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08476__A2 _03776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06487__A1 u_cpu.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10888_ _01317_ io_in[4] u_cpu.rf_ram.memory\[24\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08228__A2 _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06239__A1 _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07987__A1 _02539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05030_ u_cpu.cpu.ctrl.o_ibus_adr\[27\] _01523_ _01526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10137__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08400__A2 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07882__S _03577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05214__A2 _01704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06981_ _02957_ _03061_ _03063_ _00400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06962__A2 _03051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10287__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08720_ u_cpu.cpu.ctrl.o_ibus_adr\[30\] _04173_ _04175_ u_cpu.cpu.ctrl.o_ibus_adr\[31\]
+ _04190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05932_ _02321_ u_cpu.rf_ram.rdata\[1\] _02412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08164__A1 _03761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08651_ _03553_ _04145_ _04152_ _00982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05863_ _02341_ _02338_ _02342_ _02345_ _02346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_54_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06714__A2 _02904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07602_ _03343_ _03412_ _03413_ _00671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08582_ u_arbiter.i_wb_cpu_dbus_adr\[12\] u_arbiter.i_wb_cpu_dbus_adr\[11\] _02445_
+ _04113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_26_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05794_ _01541_ _02278_ _02279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07533_ u_cpu.rf_ram.memory\[127\]\[2\] _03372_ _03375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08467__A2 _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07464_ u_cpu.rf_ram.memory\[130\]\[7\] _03325_ _03333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06415_ u_cpu.rf_ram.memory\[47\]\[3\] _02729_ _02733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09203_ u_cpu.rf_ram.memory\[84\]\[3\] _04470_ _04477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08219__A2 _03798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07395_ _03294_ _03295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09416__A1 _04484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09134_ _04294_ _04429_ _04436_ _01181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06346_ u_cpu.rf_ram.memory\[51\]\[6\] _02686_ _02693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07978__A1 _03547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09065_ _02626_ _02727_ _04398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06277_ u_cpu.rf_ram.memory\[46\]\[1\] _02651_ _02653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08016_ _03650_ _03651_ _03655_ _00844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05228_ u_cpu.rf_ram.memory\[56\]\[1\] u_cpu.rf_ram.memory\[57\]\[1\] u_cpu.rf_ram.memory\[58\]\[1\]
+ u_cpu.rf_ram.memory\[59\]\[1\] _01602_ _01579_ _01719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06650__A1 _02742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08778__I0 _02596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05159_ _01541_ _01650_ _01651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05205__A2 _01695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09967_ _00421_ io_in[4] u_cpu.rf_ram.memory\[53\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05309__C _01426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06953__A2 _03041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09922__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08918_ _04296_ _04309_ _04317_ _01084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09898_ _00352_ io_in[4] u_cpu.rf_ram.memory\[60\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06201__S _02603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08849_ u_cpu.rf_ram.memory\[97\]\[4\] _04271_ _04276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06705__A2 _02904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10811_ _01240_ io_in[4] u_cpu.rf_ram.memory\[110\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08458__A2 _02305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06469__A1 u_arbiter.i_wb_cpu_ack vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10742_ _01171_ io_in[4] u_cpu.rf_ram.memory\[106\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07130__A2 _03139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05141__A1 _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10673_ _01102_ io_in[4] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05692__A2 _02177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07969__A1 _02561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08091__B1 _03654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05444__A2 _01932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08394__A1 _03965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07197__A2 _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06944__A2 _03041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10107_ _00553_ io_in[4] u_cpu.rf_ram.memory\[49\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11087_ _11087_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_49_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08146__A1 _01436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10038_ _00484_ io_in[4] u_cpu.rf_ram.memory\[72\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08449__A2 _03798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07121__A2 _03139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06200_ _02606_ _00076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05683__A2 _02168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06880__A1 _02963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07180_ _03175_ _03176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_129_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06131_ u_cpu.rf_ram.memory\[18\]\[6\] _02551_ _02558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09377__B _04568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06632__A1 _02742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06062_ u_cpu.rf_ram.memory\[82\]\[6\] _02477_ _02513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05013_ u_arbiter.i_wb_cpu_dbus_adr\[23\] _01442_ _01514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09945__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07188__A2 _03176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05196__I _01668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09821_ _00275_ io_in[4] u_cpu.rf_ram.memory\[6\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10922__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06935__A2 _03031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05294__S1 _01557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09752_ _00206_ io_in[4] u_cpu.rf_ram.memory\[17\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06964_ u_cpu.rf_ram.memory\[56\]\[2\] _03051_ _03054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08137__A1 _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08703_ _04181_ _01005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_55_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05915_ _01374_ _02391_ _02396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09683_ _00137_ io_in[4] u_cpu.rf_ram.memory\[51\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06895_ u_cpu.rf_ram.memory\[19\]\[3\] _03012_ _03016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06699__A1 _02561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05846_ _02305_ _02308_ _02329_ _00021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08634_ _04139_ _04142_ _04143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07360__A2 _03275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05777_ _01594_ _02261_ _01564_ _02262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08565_ _04104_ _00944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07516_ _03349_ _03362_ _03365_ _00633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08496_ u_cpu.cpu.immdec.imm19_12_20\[6\] _04016_ _04058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07112__A2 _03129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10302__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07447_ _03173_ _03315_ _03323_ _00606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08860__A2 _04282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06691__S _02894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07378_ u_cpu.rf_ram.memory\[134\]\[0\] _03285_ _03286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09117_ u_cpu.rf_ram.memory\[106\]\[7\] _04419_ _04427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06329_ _02464_ _02601_ _02682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10452__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09048_ _04388_ _04389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05977__A3 _02438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11010_ _11010_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__08376__A1 _01437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07179__A2 _02695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05809__S0 _01687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06926__A2 _03031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05285__S1 _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09242__S _04496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07351__A2 _03265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09818__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08300__A1 _03549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07103__A2 _03129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10725_ _01154_ io_in[4] u_cpu.rf_ram.memory\[79\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05114__A1 _01601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06162__I0 _02573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08851__A2 _04271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06862__A1 _02963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05665__A2 _02150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08880__I _02516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10656_ _01085_ io_in[4] u_cpu.cpu.bufreg.i_sh_signed vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08064__B1 _03678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09968__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10587_ _01017_ io_in[4] u_cpu.rf_ram.memory\[109\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05417__A2 _01877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06614__A1 _02742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04913__I _01434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10945__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06090__A2 _02530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08367__A1 _03810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04928__A1 _01437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05276__S1 _01549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07590__A2 _03402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05700_ _01422_ _02176_ _02185_ _02186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_3_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06680_ _02754_ _02884_ _02892_ _00270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07342__A2 _03265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10325__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05631_ _01539_ _02108_ _02117_ _02118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__08390__I1 u_arbiter.i_wb_cpu_rdt\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08276__B _03866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08350_ _03742_ _03768_ _03927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_17_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05562_ u_cpu.rf_ram.memory\[0\]\[5\] u_cpu.rf_ram.memory\[1\]\[5\] u_cpu.rf_ram.memory\[2\]\[5\]
+ u_cpu.rf_ram.memory\[3\]\[5\] _01556_ _01557_ _02049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_51_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09095__A2 _04409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07301_ _03171_ _03235_ _03242_ _00541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08281_ _03825_ _03870_ _03871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05493_ _01601_ _01980_ _01605_ _01981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08842__A2 _04271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10475__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07232_ _03173_ _03196_ _03204_ _00510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08055__B1 _03678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07163_ _03163_ _03159_ _03164_ _00481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05408__A2 _01896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06114_ _02512_ _02541_ _02548_ _00048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07094_ u_cpu.rf_ram.memory\[142\]\[5\] _03119_ _03125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06045_ _02477_ _02497_ _02498_ _00029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08358__A1 _03741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08358__B2 _03756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09804_ _00258_ io_in[4] u_cpu.rf_ram.memory\[76\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07030__A1 _02561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05267__S1 _01652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04919__A1 _01429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07996_ _03547_ _03636_ _03640_ _00839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07581__A2 _02821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09735_ _00189_ io_in[4] u_cpu.raddr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05592__A1 _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06947_ _02959_ _03041_ _03044_ _00385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09666_ _00120_ io_in[4] u_cpu.rf_ram.memory\[45\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06878_ _02961_ _03002_ _03006_ _00354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07333__A2 _03255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08617_ u_arbiter.i_wb_cpu_dbus_adr\[29\] u_arbiter.i_wb_cpu_dbus_adr\[28\] _04115_
+ _04131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05344__A1 _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05829_ u_cpu.cpu.decode.opcode\[0\] _02313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09597_ _00051_ io_in[4] u_cpu.rf_ram.memory\[18\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05895__A2 u_cpu.cpu.ctrl.i_iscomp vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10818__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08548_ u_cpu.rf_ram.memory\[31\]\[1\] _04094_ _04096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09086__A2 _04409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07097__A1 _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08479_ _03828_ _03818_ _03788_ _04042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10510_ _00943_ io_in[4] u_cpu.cpu.alu.cmp_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06844__A1 _02963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07892__I0 _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10441_ _00874_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08046__B1 _03676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10372_ _00805_ io_in[4] u_cpu.rf_ram.memory\[112\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08141__S _01434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05992__C _01373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09010__A2 _04359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07021__A1 _02961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07572__A2 _03392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10348__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09640__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08521__A1 _03798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07324__A2 _03255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05335__A1 _01636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10498__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05513__B _01626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05886__A2 _01369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09077__A2 _04399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09790__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10708_ _01137_ io_in[4] u_cpu.rf_ram.memory\[104\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10639_ _01068_ io_in[4] u_cpu.rf_ram.memory\[94\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06063__A2 _02512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05497__S1 _01616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05810__A2 _02294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09001__A2 _04359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07012__A1 _02524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07850_ _03543_ _03558_ _03560_ _00773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07563__A2 _02821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07890__S _03577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06801_ u_cpu.rf_ram.memory\[29\]\[3\] _02955_ _02962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07781_ u_cpu.rf_ram.memory\[35\]\[7\] _03510_ _03518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04993_ u_cpu.cpu.ctrl.o_ibus_adr\[19\] _01495_ _01498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_83_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09520_ u_cpu.rf_ram.memory\[100\]\[6\] _04654_ _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06732_ _02752_ _02914_ _02921_ _00293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08512__A1 _03741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07315__A2 _03245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08512__B2 _03791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05326__A1 _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09451_ u_cpu.rf_ram.memory\[25\]\[7\] _04615_ _04623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06663_ _02626_ _02706_ _02883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05614_ _01398_ _02100_ _02101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08402_ _03973_ _03851_ _03826_ _03974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_80_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09382_ _04580_ _04581_ _04582_ _02349_ _01283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06594_ _02738_ _02844_ _02845_ _00231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09068__A2 _04399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08333_ _01380_ _03740_ _03913_ _00903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05545_ u_cpu.rf_ram.memory\[136\]\[4\] u_cpu.rf_ram.memory\[137\]\[4\] u_cpu.rf_ram.memory\[138\]\[4\]
+ u_cpu.rf_ram.memory\[139\]\[4\] _01680_ _01681_ _02033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_20_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08815__A2 _03769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08264_ _01381_ _03740_ _03855_ _00892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06826__A1 _02963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05476_ _01957_ _01959_ _01961_ _01963_ _01568_ _01964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_137_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07215_ _02626_ _02893_ _03195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08195_ _02383_ _03740_ _03794_ _00884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07146_ _03153_ _00475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_3_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07251__A1 _02577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07077_ _03115_ _00444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05488__S1 _01548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06028_ _02478_ u_cpu.rf_ram_if.wdata1_r\[1\] _02484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07003__A1 _02961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09663__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07554__A2 _03382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07979_ u_cpu.rf_ram.memory\[116\]\[4\] _03626_ _03631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09718_ _00172_ io_in[4] u_cpu.rf_ram.memory\[50\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10990_ _10990_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__10640__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08503__A1 _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07306__A2 _03245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08628__C _02773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09649_ _00103_ io_in[4] u_cpu.rf_ram.memory\[42\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05317__A1 _01601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05333__B _01416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09059__A2 _04389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10790__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07490__A1 _03347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10020__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10424_ _00857_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09231__A2 _04487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06045__A2 _02497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07242__A1 _03165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05479__S1 _01580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10355_ _00788_ io_in[4] u_cpu.rf_ram.memory\[8\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07793__A2 _03520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08990__A1 _04294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10286_ _00719_ io_in[4] u_cpu.rf_ram.memory\[90\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10170__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xu_scanchain_local.scan_flop\[12\] u_arbiter.i_wb_cpu_rdt\[9\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[6\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_78_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07545__A2 _02821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05100__S0 _01590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09298__A2 _04526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05308__A1 _01542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05330_ u_cpu.rf_ram.memory\[108\]\[2\] u_cpu.rf_ram.memory\[109\]\[2\] u_cpu.rf_ram.memory\[110\]\[2\]
+ u_cpu.rf_ram.memory\[111\]\[2\] _01598_ _01620_ _01820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06808__A1 _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09470__A2 _04625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06284__A2 _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05261_ u_cpu.rf_ram.memory\[92\]\[1\] u_cpu.rf_ram.memory\[93\]\[1\] u_cpu.rf_ram.memory\[94\]\[1\]
+ u_cpu.rf_ram.memory\[95\]\[1\] _01610_ _01611_ _01752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_30_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07000_ u_cpu.rf_ram.memory\[54\]\[2\] _03071_ _03074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05192_ _01667_ _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08025__A3 u_arbiter.i_wb_cpu_dbus_dat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09222__A2 _04487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10513__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07233__A1 _02727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07684__I _02783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09686__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08951_ u_arbiter.i_wb_cpu_rdt\[20\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[4\]
+ _04331_ _04336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_124_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07902_ _03588_ _00797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08882_ _04296_ _04282_ _04297_ _01068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10663__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08733__A1 _03539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07536__A2 _03372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07833_ _02501_ _03549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05137__C _01628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07764_ _03359_ _03500_ _03508_ _00739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04976_ _01483_ _01485_ u_arbiter.o_wb_cpu_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09503_ _04482_ _04644_ _04651_ _01335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06715_ u_cpu.rf_ram.memory\[68\]\[7\] _02904_ _02912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07695_ _03343_ _03465_ _03466_ _00711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09434_ _04484_ _04605_ _04613_ _01304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06646_ _02873_ _02874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_24_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09365_ _01385_ u_cpu.cpu.genblk3.csr.mcause3_0\[1\] _04570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06577_ u_cpu.rf_ram.memory\[129\]\[1\] _02834_ _02836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10043__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08316_ _03785_ _03896_ _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05528_ _01645_ _02015_ _01648_ _02016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05158__S0 _01590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09296_ u_cpu.rf_ram.memory\[86\]\[3\] _04526_ _04530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09461__A2 _04625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06275__A2 _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08247_ _02332_ _03740_ _03840_ _00890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05459_ u_cpu.rf_ram.memory\[140\]\[3\] u_cpu.rf_ram.memory\[141\]\[3\] u_cpu.rf_ram.memory\[142\]\[3\]
+ u_cpu.rf_ram.memory\[143\]\[3\] _01680_ _01681_ _01948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_119_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10193__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08178_ _02765_ u_arbiter.i_wb_cpu_rdt\[15\] _03777_ _03778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_u_scanchain_local.scan_flop\[10\]_D u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09213__A2 _04470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06027__A2 _02482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07224__A1 _03165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07129_ _02963_ _03139_ _03144_ _00467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07775__A2 _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10140_ _00586_ io_in[4] u_cpu.rf_ram.memory\[133\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05786__A1 _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05330__S0 _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10071_ _00517_ io_in[4] u_cpu.rf_ram.memory\[143\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07527__A2 _02821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[14\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06003__I u_cpu.rf_ram_if.genblk1.wtrig0_r vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05633__S1 _01681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10973_ _10973_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_71_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09250__S _04496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05998__B _02332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09452__A2 _04615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10536__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06266__A2 _02641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07463__A1 _03171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08660__B1 _04157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[8\]_D u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09204__A2 _04470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07215__A1 _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10407_ _00840_ io_in[4] u_cpu.rf_ram.memory\[33\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10686__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04921__I _01442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10338_ _00771_ io_in[4] u_cpu.rf_ram.memory\[120\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05321__S0 _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05777__A1 _01594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05238__B _01626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10269_ _00702_ io_in[4] u_cpu.rf_ram.memory\[36\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07518__A2 _03362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08191__A2 _03755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05624__S1 _01652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09140__A1 _04280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10066__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06500_ u_cpu.rf_ram.memory\[16\]\[0\] _02791_ _02792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07480_ _03341_ _00621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06431_ u_cpu.rf_ram.memory\[50\]\[1\] _02740_ _02743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06362_ _02502_ _02697_ _02702_ _00142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09150_ _04292_ _04439_ _04445_ _01188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09443__A2 _04615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08101_ _03715_ _03716_ _00868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05313_ _01594_ _01802_ _01564_ _01803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06257__A2 _02641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06293_ _02661_ _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09081_ u_cpu.rf_ram.memory\[79\]\[7\] _04399_ _04407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05244_ u_cpu.rf_ram.memory\[104\]\[1\] u_cpu.rf_ram.memory\[105\]\[1\] u_cpu.rf_ram.memory\[106\]\[1\]
+ u_cpu.rf_ram.memory\[107\]\[1\] _01615_ _01616_ _01735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_107_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08032_ _03653_ _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05560__S0 _01546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07206__A1 _03165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08254__I0 u_arbiter.i_wb_cpu_rdt\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05175_ _01540_ _01667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07757__A2 _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[37\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09983_ _00437_ io_in[4] u_cpu.rf_ram.memory\[9\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05768__A1 _01421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05312__S0 _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05148__B _01626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08934_ u_cpu.rf_ram.memory\[28\]\[4\] _04322_ _04327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07509__A2 _02832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08865_ _02491_ _04286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__04991__A2 _01442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10409__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07816_ _03357_ _03530_ _03537_ _00762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05615__S1 _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08796_ u_cpu.rf_ram.memory\[93\]\[6\] _04227_ _04234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07747_ _02475_ _02671_ _03499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04959_ u_cpu.cpu.ctrl.o_ibus_adr\[10\] _01471_ _01472_ _01473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05940__A1 _02320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09701__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07678_ u_cpu.cpu.mem_bytecnt\[0\] _03454_ _03455_ _00705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_41_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10559__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09417_ _02528_ _02638_ _04604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06629_ u_cpu.rf_ram.memory\[74\]\[0\] _02864_ _02865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09348_ u_cpu.rf_ram.memory\[88\]\[2\] _04556_ _04559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09851__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09434__A2 _04605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06248__A2 _02628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07445__A1 _03171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09279_ _04476_ _04516_ _04520_ _01242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07996__A2 _03636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05551__S0 _01687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09198__A1 _04472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05303__S0 _01578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06420__A2 _02729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10123_ _00569_ io_in[4] u_cpu.rf_ram.memory\[135\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10054_ _00500_ io_in[4] u_cpu.rf_ram.memory\[71\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[5\] u_arbiter.i_wb_cpu_rdt\[2\] io_in[3] u_arbiter.i_wb_cpu_dbus_sel\[3\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_75_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10089__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07920__A2 _03596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09122__A1 _04280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10956_ u_cpu.cpu.o_wen1 io_in[4] u_cpu.rf_ram_if.wen1_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06487__A2 _01385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10887_ _01316_ io_in[4] u_cpu.rf_ram.memory\[24\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09425__A2 _04605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06239__A2 _02628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07987__A2 _02639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05998__A1 _02431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06411__A2 _02729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06980_ u_cpu.rf_ram.memory\[55\]\[1\] _03061_ _03063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05931_ _02411_ u_cpu.cpu.o_wdata0 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_79_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04973__A2 _01443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09724__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08164__A2 _03762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09361__A1 _02305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08650_ u_cpu.rf_ram.memory\[30\]\[6\] _04145_ _04152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05862_ _02305_ _02344_ _02345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07601_ u_cpu.rf_ram.memory\[123\]\[0\] _03412_ _03413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05415__C _01628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08581_ _04112_ _00952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_81_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05793_ u_cpu.rf_ram.memory\[80\]\[7\] u_cpu.rf_ram.memory\[81\]\[7\] u_cpu.rf_ram.memory\[82\]\[7\]
+ u_cpu.rf_ram.memory\[83\]\[7\] _01590_ _01591_ _02278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10701__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07532_ _03347_ _03372_ _03374_ _00640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09874__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06478__A2 _02773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07463_ _03171_ _03325_ _03332_ _00613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09202_ _02496_ _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06414_ _02492_ _02729_ _02732_ _00164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10851__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07394_ _02524_ _02832_ _03294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05781__S0 _01646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09416__A2 _04595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09133_ u_cpu.rf_ram.memory\[107\]\[6\] _04429_ _04436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07427__A1 _03171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06345_ _02507_ _02686_ _02692_ _00135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07978__A2 _03626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09064_ _04296_ _04389_ _04397_ _01150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06276_ _02482_ _02651_ _02652_ _00106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08015_ u_arbiter.i_wb_cpu_rdt\[0\] _03653_ _03654_ u_arbiter.i_wb_cpu_dbus_dat\[0\]
+ _03655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05227_ _01597_ _01717_ _01718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06650__A2 _02874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08927__A1 _04280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05158_ u_cpu.rf_ram.memory\[112\]\[0\] u_cpu.rf_ram.memory\[113\]\[0\] u_cpu.rf_ram.memory\[114\]\[0\]
+ u_cpu.rf_ram.memory\[115\]\[0\] _01590_ _01591_ _01650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_116_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06402__A2 _02718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10231__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06689__S _02894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09966_ _00420_ io_in[4] u_cpu.rf_ram.memory\[53\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05089_ u_cpu.rf_ram.memory\[16\]\[0\] u_cpu.rf_ram.memory\[17\]\[0\] u_cpu.rf_ram.memory\[18\]\[0\]
+ u_cpu.rf_ram.memory\[19\]\[0\] _01578_ _01580_ _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_58_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08917_ u_cpu.rf_ram.memory\[96\]\[7\] _04309_ _04317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04964__A2 _01457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09897_ _00351_ io_in[4] u_cpu.rf_ram.memory\[60\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08848_ _03547_ _04271_ _04275_ _01056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05606__B _01648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10381__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05913__A1 _02311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08779_ _04224_ _01038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_45_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09104__A1 _04280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10810_ _01239_ io_in[4] u_cpu.rf_ram.memory\[110\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08458__A3 _03798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10741_ _01170_ io_in[4] u_cpu.rf_ram.memory\[106\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07666__A1 _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06469__A2 _01431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05141__A2 _01632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10672_ _01101_ io_in[4] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05772__S0 _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09407__A2 _04595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07969__A2 _02821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08091__A1 u_arbiter.i_wb_cpu_rdt\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08144__S _01434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06641__A2 _02864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08918__A1 _04296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09747__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[42\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10106_ _00552_ io_in[4] u_cpu.rf_ram.memory\[49\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11086_ _11086_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_110_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04955__A2 _01443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10724__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10037_ _00483_ io_in[4] u_cpu.rf_ram.memory\[72\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06157__A1 u_cpu.cpu.immdec.imm11_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09897__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[57\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10874__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10939_ u_cpu.rf_ram_if.wdata0_r\[6\] io_in[4] u_cpu.rf_ram_if.wdata0_r\[5\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05763__S0 _01619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10104__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07409__A1 _03171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06880__A2 _03002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06130_ _02507_ _02551_ _02557_ _00055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05515__S0 _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06061_ _02511_ _02512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06632__A2 _02864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10254__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05012_ _01507_ _01512_ _01513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09820_ _00274_ io_in[4] u_cpu.rf_ram.memory\[6\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09751_ _00205_ io_in[4] u_cpu.rf_ram.memory\[17\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06963_ _02957_ _03051_ _03053_ _00392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08137__A2 _03731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08702_ u_cpu.cpu.ctrl.o_ibus_adr\[21\] _04173_ _04175_ u_cpu.cpu.ctrl.o_ibus_adr\[22\]
+ _04181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_104_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05914_ u_cpu.cpu.state.o_cnt\[2\] u_cpu.cpu.mem_bytecnt\[0\] _02395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_67_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06148__A1 _02502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09682_ _00136_ io_in[4] u_cpu.rf_ram.memory\[51\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06894_ _02959_ _03012_ _03015_ _00361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08633_ _04137_ _04141_ _04142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05845_ _02305_ _02328_ _02329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06699__A2 _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08564_ u_arbiter.i_wb_cpu_dbus_adr\[3\] u_arbiter.i_wb_cpu_dbus_adr\[2\] _02445_
+ _04104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05776_ u_cpu.rf_ram.memory\[96\]\[7\] u_cpu.rf_ram.memory\[97\]\[7\] u_cpu.rf_ram.memory\[98\]\[7\]
+ u_cpu.rf_ram.memory\[99\]\[7\] _01602_ _01579_ _02261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_74_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07648__A1 _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07515_ u_cpu.rf_ram.memory\[128\]\[2\] _03362_ _03365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08495_ u_cpu.cpu.immdec.imm19_12_20\[7\] _02768_ _04057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_23_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07446_ u_cpu.rf_ram.memory\[131\]\[7\] _03315_ _03323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06320__A1 _02497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05754__S0 _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07377_ _03284_ _03285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06871__A2 _03002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08472__B _04016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09116_ _04294_ _04419_ _04426_ _01173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06328_ _02517_ _02673_ _02681_ _00129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05506__S0 _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09047_ _02682_ _04197_ _04388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07820__A1 _02810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06623__A2 _02854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06259_ u_cpu.rf_ram.memory\[42\]\[1\] _02641_ _02643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10747__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08376__A2 u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05809__S1 _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06387__A1 _02517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09949_ _00403_ io_in[4] u_cpu.rf_ram.memory\[55\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08128__A2 _03731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10897__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05850__I u_cpu.cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10127__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08300__A2 _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10724_ _01153_ io_in[4] u_cpu.rf_ram.memory\[79\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06311__A1 _02639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05114__A2 _01604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05745__S0 _01546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10655_ _01084_ io_in[4] u_cpu.rf_ram.memory\[96\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06862__A2 _02992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10277__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08064__A1 u_arbiter.i_wb_cpu_rdt\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10586_ _01016_ io_in[4] u_cpu.rf_ram.memory\[109\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xu_scanchain_local.scan_flop\[42\] u_scanchain_local.module_data_in\[41\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[4\] u_scanchain_local.clk u_scanchain_local.module_data_in\[42\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__05417__A3 _01886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06614__A2 _02854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08119__A2 _03678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11069_ _11069_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_3_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07878__A1 _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05630_ _02110_ _02112_ _02114_ _02116_ _01568_ _02117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_24_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06550__A1 _02752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05561_ _01554_ _02047_ _02048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07300_ u_cpu.rf_ram.memory\[39\]\[6\] _03235_ _03242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07888__S _03577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08280_ _03791_ _03869_ _03870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05492_ u_cpu.rf_ram.memory\[56\]\[4\] u_cpu.rf_ram.memory\[57\]\[4\] u_cpu.rf_ram.memory\[58\]\[4\]
+ u_cpu.rf_ram.memory\[59\]\[4\] _01602_ _01579_ _01980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__05736__S0 _01578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07231_ u_cpu.rf_ram.memory\[70\]\[7\] _03196_ _03204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09388__B _01429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06853__A2 _02992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09912__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08055__A1 u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07162_ u_cpu.rf_ram.memory\[72\]\[2\] _03159_ _03164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08055__B2 u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06113_ u_cpu.rf_ram.memory\[81\]\[6\] _02541_ _02548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07093_ _02963_ _03119_ _03124_ _00451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06605__A2 _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06044_ u_cpu.rf_ram.memory\[82\]\[3\] _02477_ _02498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09555__A1 _04480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08358__A2 _03786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09803_ _00257_ io_in[4] u_cpu.rf_ram.memory\[76\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_101_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07030__A2 _02684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07995_ u_cpu.rf_ram.memory\[33\]\[3\] _03636_ _03640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05041__A1 _01443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09734_ _00188_ io_in[4] u_cpu.rf_ram_if.rcnt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06946_ u_cpu.rf_ram.memory\[57\]\[2\] _03041_ _03044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09665_ _00119_ io_in[4] u_cpu.rf_ram.memory\[45\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06916__I0 _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06877_ u_cpu.rf_ram.memory\[60\]\[3\] _03002_ _03006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08530__A2 _04084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08616_ _04130_ _00969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05828_ u_cpu.cpu.immdec.imm11_7\[0\] _02312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_82_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09596_ _00050_ io_in[4] u_cpu.rf_ram.memory\[18\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08547_ _03539_ _04094_ _04095_ _00935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05759_ u_cpu.rf_ram.memory\[40\]\[7\] u_cpu.rf_ram.memory\[41\]\[7\] u_cpu.rf_ram.memory\[42\]\[7\]
+ u_cpu.rf_ram.memory\[43\]\[7\] _01545_ _01642_ _02244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_126_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08294__A1 _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07097__A2 _03119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08478_ _03756_ _03789_ _03892_ _04041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05727__S0 _01687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09592__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07429_ _03173_ _03305_ _03313_ _00598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06844__A2 _02982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08046__A1 u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10440_ _00873_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08046__B2 _02779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06207__S _02603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10371_ _00804_ io_in[4] u_cpu.rf_ram.memory\[112\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05280__A1 _01751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07021__A2 _03081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06780__A1 _02746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08521__A2 _03906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09935__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08285__A1 _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07088__A2 _03119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10707_ _01136_ io_in[4] u_cpu.rf_ram.memory\[104\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10912__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06835__A2 _02982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10638_ _01067_ io_in[4] u_cpu.rf_ram.memory\[94\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__04924__I _01442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10569_ _00999_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05271__A1 _01667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09537__A1 _04480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07012__A2 _02684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06800_ _02496_ _02961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07780_ _03357_ _03510_ _03517_ _00746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_04992_ _01443_ _01495_ _01496_ _01497_ u_arbiter.o_wb_cpu_adr\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__06771__A1 _02612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06731_ u_cpu.rf_ram.memory\[67\]\[6\] _02914_ _02921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09450_ _04482_ _04615_ _04622_ _01311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05704__B _01648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06662_ _02754_ _02874_ _02882_ _00262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10442__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05326__A2 _01815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06523__A1 _02744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08401_ _02765_ u_arbiter.i_wb_cpu_rdt\[9\] _03972_ _03973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_24_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05613_ u_cpu.rf_ram.memory\[92\]\[5\] u_cpu.rf_ram.memory\[93\]\[5\] u_cpu.rf_ram.memory\[94\]\[5\]
+ u_cpu.rf_ram.memory\[95\]\[5\] _01610_ _01611_ _02100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_91_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09381_ u_cpu.cpu.genblk3.csr.o_new_irq _04581_ _04582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05877__A3 _02325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06593_ u_cpu.rf_ram.memory\[139\]\[0\] _02844_ _02845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08332_ _03889_ _03912_ _03913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05544_ _02012_ _02031_ _01402_ _02032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08276__A1 _02343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10592__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08263_ _03816_ _03846_ _03854_ _03855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06826__A2 _02972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05475_ _01562_ _01962_ _01565_ _01963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07214_ _03173_ _03186_ _03194_ _00502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08194_ _03740_ _03793_ _03794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07145_ _02590_ u_cpu.rf_ram.memory\[13\]\[4\] _03148_ _03153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05637__I0 u_cpu.rf_ram.memory\[128\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07076_ _02593_ u_cpu.rf_ram.memory\[15\]\[5\] _03109_ _03115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07251__A2 _02625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05262__A1 _01398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06027_ _02477_ _02482_ _02483_ _00026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09808__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08200__A1 _01436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07003__A2 _03071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05014__A1 _01443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07978_ _03547_ _03626_ _03630_ _00831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06697__S _02894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06762__A1 _02746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09717_ _00171_ io_in[4] u_cpu.rf_ram.memory\[50\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06929_ _02959_ _03031_ _03034_ _00377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09958__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08503__A2 _04059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09648_ _00102_ io_in[4] u_cpu.rf_ram.memory\[42\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05317__A2 _01806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09579_ _00033_ io_in[4] u_cpu.rf_ram.memory\[82\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10935__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08267__A1 _03831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06817__A2 _02972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08019__A1 _03648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07490__A2 _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10423_ _00856_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09248__S _04496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10354_ _00787_ io_in[4] u_cpu.rf_ram.memory\[121\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07242__A2 _03206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10315__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09519__A1 _04480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08990__A2 _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10285_ _00718_ io_in[4] u_cpu.rf_ram.memory\[91\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08742__A2 _04199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10465__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05100__S1 _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06753__A1 _02539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06505__A1 _02744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05308__A2 _01797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08258__A1 _03773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06808__A2 _02955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05260_ _01422_ _01741_ _01750_ _01751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_128_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05191_ _01399_ _01682_ _01683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07233__A2 _02832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08430__A1 _02765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08981__A2 _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08950_ _04335_ _01098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10808__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07901_ _02581_ u_cpu.rf_ram.memory\[11\]\[1\] _03586_ _03588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08881_ u_cpu.rf_ram.memory\[94\]\[7\] _04282_ _04297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07832_ _03547_ _03541_ _03548_ _00767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08733__A2 _04199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06744__A1 _02746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07763_ u_cpu.rf_ram.memory\[92\]\[7\] _03500_ _03508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04975_ u_cpu.cpu.ctrl.o_ibus_adr\[14\] _01481_ _01484_ _01485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09502_ u_cpu.rf_ram.memory\[98\]\[6\] _04644_ _04651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06714_ _02752_ _02904_ _02911_ _00285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05434__B _01654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08497__A1 _04016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07694_ u_cpu.rf_ram.memory\[91\]\[0\] _03465_ _03466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09433_ u_cpu.rf_ram.memory\[26\]\[7\] _04605_ _04613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06645_ _02626_ _02671_ _02873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09364_ u_cpu.cpu.genblk3.csr.o_new_irq _01392_ _04569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06576_ _02738_ _02834_ _02835_ _00223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07141__S _03148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08315_ _03776_ _03768_ _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05527_ u_cpu.rf_ram.memory\[88\]\[4\] u_cpu.rf_ram.memory\[89\]\[4\] u_cpu.rf_ram.memory\[90\]\[4\]
+ u_cpu.rf_ram.memory\[91\]\[4\] _01646_ _01603_ _02015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09295_ _04474_ _04526_ _04529_ _01249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05158__S1 _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08246_ _03811_ _03802_ _03839_ _02768_ _03840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_36_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05458_ _01399_ _01946_ _01947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10338__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08177_ _01435_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\] _03777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_119_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05389_ u_cpu.rf_ram.memory\[20\]\[3\] u_cpu.rf_ram.memory\[21\]\[3\] u_cpu.rf_ram.memory\[22\]\[3\]
+ u_cpu.rf_ram.memory\[23\]\[3\] _01572_ _01574_ _01878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_118_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09630__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07128_ u_cpu.rf_ram.memory\[140\]\[4\] _03139_ _03144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07224__A2 _03196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08421__A1 _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08421__B2 _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07059_ _02593_ u_cpu.rf_ram.memory\[9\]\[5\] _03100_ _03106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10488__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05330__S1 _01620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06983__A1 _02959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10070_ _00516_ io_in[4] u_cpu.rf_ram.memory\[143\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09780__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06735__A1 _02469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05094__S0 _01578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10972_ _10972_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_16_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07160__A1 _03161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07051__S _03100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08660__A1 u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07463__A2 _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10406_ _00839_ io_in[4] u_cpu.rf_ram.memory\[33\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07215__A2 _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10337_ _00770_ io_in[4] u_cpu.rf_ram.memory\[120\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05777__A2 _02261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05321__S1 _01616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10268_ _00701_ io_in[4] u_cpu.rf_ram.memory\[36\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10199_ _00645_ io_in[4] u_cpu.rf_ram.memory\[127\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06726__A1 _02746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05254__B _01648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08479__A1 _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09140__A2 _04439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06430_ _02486_ _02742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08284__C _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06361_ u_cpu.rf_ram.memory\[41\]\[4\] _02697_ _02702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08100__B1 _03676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08100_ u_arbiter.i_wb_cpu_dbus_dat\[24\] _03654_ _03676_ u_arbiter.i_wb_cpu_dbus_dat\[25\]
+ _03716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07896__S _03577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05312_ u_cpu.rf_ram.memory\[48\]\[2\] u_cpu.rf_ram.memory\[49\]\[2\] u_cpu.rf_ram.memory\[50\]\[2\]
+ u_cpu.rf_ram.memory\[51\]\[2\] _01544_ _01548_ _01802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09653__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09080_ _04294_ _04399_ _04406_ _01157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06292_ _02639_ _02660_ _02661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07454__A2 _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08651__A1 _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08031_ u_arbiter.i_wb_cpu_rdt\[3\] _03668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05243_ _01597_ _01733_ _01734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05560__S1 _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10630__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07206__A2 _03186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08403__A1 _03812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05174_ _01659_ _01661_ _01663_ _01665_ _01426_ _01666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__08254__I1 u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09982_ _00436_ io_in[4] u_cpu.rf_ram.memory\[9\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06965__A1 _02959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05312__S1 _01548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08933_ _04288_ _04322_ _04326_ _01090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10780__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08706__A2 _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08864_ _04284_ _04282_ _04285_ _01062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06717__A1 _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07815_ u_cpu.rf_ram.memory\[117\]\[6\] _03530_ _03537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08795_ _03551_ _04227_ _04233_ _01045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10010__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07746_ _01428_ _03451_ _03498_ _00731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_04958_ u_cpu.cpu.ctrl.o_ibus_adr\[10\] _01471_ _01442_ _01472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_84_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09131__A2 _04429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07677_ u_cpu.cpu.mem_bytecnt\[0\] _03454_ _01429_ _03455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_04889_ _01407_ _01414_ _01415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_13_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09416_ _04484_ _04595_ _04603_ _01296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06628_ _02863_ _02864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08890__A1 _04286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10160__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09347_ _04472_ _04556_ _04558_ _01272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05611__C _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06559_ _02742_ _02823_ _02825_ _00216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09278_ u_cpu.rf_ram.memory\[110\]\[3\] _04516_ _04520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07445__A2 _03315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05456__A1 _01925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08229_ _03771_ _03813_ _03816_ _03757_ _03824_ _00888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_126_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05551__S1 _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09198__A2 _04470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05303__S1 _01580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10122_ _00568_ io_in[4] u_cpu.rf_ram.memory\[135\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10053_ _00499_ io_in[4] u_cpu.rf_ram.memory\[71\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06708__A1 _02746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07381__A1 _03161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05074__B _01565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09122__A2 _04429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10955_ u_cpu.cpu.o_wen0 io_in[4] u_cpu.rf_ram_if.wen0_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10503__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07133__A1 _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09676__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06487__A3 _02433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10886_ _01315_ io_in[4] u_cpu.rf_ram.memory\[24\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10653__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08633__A1 _04137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07436__A2 _03315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08605__S _04115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05447__A1 _01667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09189__A2 _04459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05249__B _01626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08936__A2 _04322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06947__A1 _02959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05930_ _01386_ _02408_ _02410_ _02411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10033__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08164__A3 _03763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09361__A2 _02344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05861_ _02343_ u_cpu.cpu.decode.co_ebreak _01411_ _02344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_113_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07600_ _03411_ _03412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08580_ u_arbiter.i_wb_cpu_dbus_adr\[11\] u_arbiter.i_wb_cpu_dbus_adr\[10\] _02445_
+ _04112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05792_ _01645_ _02276_ _01648_ _02277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07531_ u_cpu.rf_ram.memory\[127\]\[1\] _03372_ _03374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09113__A2 _04419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10183__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08172__I0 u_arbiter.i_wb_cpu_rdt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07462_ u_cpu.rf_ram.memory\[130\]\[6\] _03325_ _03332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07675__A2 u_cpu.cpu.state.o_cnt_r\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09201_ _04474_ _04470_ _04475_ _01209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06413_ u_cpu.rf_ram.memory\[47\]\[2\] _02729_ _02732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07393_ _03173_ _03285_ _03293_ _00582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05781__S1 _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09132_ _04292_ _04429_ _04435_ _01180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06344_ u_cpu.rf_ram.memory\[51\]\[5\] _02686_ _02692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08624__A1 u_cpu.cpu.bufreg.i_sh_signed vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07427__A2 _03305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05438__A1 _01398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09063_ u_cpu.rf_ram.memory\[99\]\[7\] _04389_ _04397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06275_ u_cpu.rf_ram.memory\[46\]\[0\] _02651_ _02652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08014_ _03653_ _03648_ _03654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05226_ u_cpu.rf_ram.memory\[60\]\[1\] u_cpu.rf_ram.memory\[61\]\[1\] u_cpu.rf_ram.memory\[62\]\[1\]
+ u_cpu.rf_ram.memory\[63\]\[1\] _01598_ _01573_ _01717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_118_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08927__A2 _04322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05157_ _01645_ _01647_ _01648_ _01649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09965_ _00419_ io_in[4] u_cpu.rf_ram.memory\[53\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05088_ _01579_ _01580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05610__A1 _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08916_ _04294_ _04309_ _04316_ _01083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09896_ _00350_ io_in[4] u_cpu.rf_ram.memory\[61\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09352__A2 _04556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08847_ u_cpu.rf_ram.memory\[97\]\[3\] _04271_ _04275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10526__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[11\]_SI u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07363__A1 _03161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09699__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08778_ _02596_ u_cpu.rf_ram.memory\[2\]\[6\] _04217_ _04224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_57_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09104__A2 _04419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07729_ u_cpu.cpu.state.genblk1.misalign_trap_sync_r _03458_ _03485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07115__A1 _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08163__I0 u_arbiter.i_wb_cpu_rdt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10740_ _01169_ io_in[4] u_cpu.rf_ram.memory\[106\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10676__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07666__A2 _03442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10671_ _01100_ io_in[4] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05772__S1 _01616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07418__A2 _03305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08091__A2 _03653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08918__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10056__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09040__A1 _04290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06929__A1 _02959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05601__A1 _01594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10105_ _00551_ io_in[4] u_cpu.rf_ram.memory\[49\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11085_ _11085_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_95_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10036_ _00482_ io_in[4] u_cpu.rf_ram.memory\[72\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05532__B _01654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08854__A1 _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07657__A2 _03442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[27\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10938_ u_cpu.rf_ram_if.wdata0_r\[5\] io_in[4] u_cpu.rf_ram_if.wdata0_r\[4\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07901__I0 _02581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10869_ _01298_ io_in[4] u_cpu.rf_ram.memory\[26\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05763__S1 _01620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07409__A2 _03295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08082__A2 _03683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05515__S1 _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06093__A1 _02507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06060_ _02510_ _02511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05011_ u_cpu.cpu.ctrl.o_ibus_adr\[23\] u_cpu.cpu.ctrl.o_ibus_adr\[22\] _01512_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05840__A1 _02320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08909__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10549__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06396__A2 _02718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06962_ u_cpu.rf_ram.memory\[56\]\[1\] _03051_ _03053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09750_ _00204_ io_in[4] u_cpu.rf_ram.memory\[17\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09841__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09334__A2 _04546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05913_ _02311_ _02392_ _02393_ _02394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08701_ _04180_ _01004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_39_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09681_ _00135_ io_in[4] u_cpu.rf_ram.memory\[51\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05426__C _01628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06893_ u_cpu.rf_ram.memory\[19\]\[2\] _03012_ _03015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06148__A2 _02563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07345__A1 _03161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08632_ u_arbiter.i_wb_cpu_dbus_adr\[2\] _02448_ _04141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10699__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05844_ _02310_ _02326_ _02327_ _02328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08563_ _02433_ _03494_ _04103_ _00943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09098__A1 _04294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05775_ _01636_ _02259_ _02260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09991__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07514_ _03347_ _03362_ _03364_ _00632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07648__A2 _03432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08494_ _03782_ _04050_ _04052_ _04055_ _03797_ _04056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_50_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07445_ _03171_ _03315_ _03322_ _00605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06320__A2 _02673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05754__S1 _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07376_ _02832_ _02893_ _03284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09115_ u_cpu.rf_ram.memory\[106\]\[6\] _04419_ _04426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06327_ u_cpu.rf_ram.memory\[44\]\[7\] _02673_ _02681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10079__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09270__A1 _02625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05506__S1 _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09046_ _04296_ _04379_ _04387_ _01142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06258_ _02482_ _02641_ _02642_ _00098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07820__A2 _02821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05209_ _01554_ _01699_ _01700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05831__A1 _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09022__A1 _04290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06189_ _02598_ _02599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07584__A1 _03343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06387__A2 _02708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09948_ _00402_ io_in[4] u_cpu.rf_ram.memory\[55\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09879_ _00333_ io_in[4] u_cpu.rf_ram.memory\[63\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06139__A2 _02563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05898__A1 u_arbiter.i_wb_cpu_ibus_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05352__B _01648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07639__A2 _03432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08836__A1 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10723_ _01152_ io_in[4] u_cpu.rf_ram.memory\[79\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06311__A2 _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05745__S1 _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10654_ _01083_ io_in[4] u_cpu.rf_ram.memory\[96\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08155__S _01435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09714__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09261__A1 _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08064__A2 _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10585_ _01015_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07811__A2 _03530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[35\] u_scanchain_local.module_data_in\[34\] io_in[3]
+ u_arbiter.i_wb_cpu_dbus_dat\[29\] u_scanchain_local.clk u_scanchain_local.module_data_in\[35\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_123_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09864__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08611__I1 u_arbiter.i_wb_cpu_dbus_adr\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06378__A2 _02708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10841__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09316__A2 _04536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11068_ _11068_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_23_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07327__A1 _03161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10019_ _00465_ io_in[4] u_cpu.rf_ram.memory\[140\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05338__B1 _01825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07878__A2 _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05433__S0 _01623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06550__A2 _02812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05560_ u_cpu.rf_ram.memory\[4\]\[5\] u_cpu.rf_ram.memory\[5\]\[5\] u_cpu.rf_ram.memory\[6\]\[5\]
+ u_cpu.rf_ram.memory\[7\]\[5\] _01546_ _01550_ _02047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08827__A1 _03778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08827__B2 _03742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06689__I0 _02587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05491_ _01597_ _01978_ _01979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06302__A2 _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05736__S1 _01580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10221__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07230_ _03171_ _03196_ _03203_ _00509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07161_ _02491_ _03163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09252__A1 _02475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08055__A2 _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06112_ _02507_ _02541_ _02547_ _00047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07092_ u_cpu.rf_ram.memory\[142\]\[4\] _03119_ _03124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10371__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06043_ _02496_ _02497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09004__A1 _04290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09555__A2 _04674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07566__A1 _03343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09802_ _00256_ io_in[4] u_cpu.rf_ram.memory\[76\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07994_ _03545_ _03636_ _03639_ _00838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09733_ _00187_ io_in[4] u_cpu.rf_ram_if.rcnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06945_ _02957_ _03041_ _03043_ _00384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05592__A3 _02078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07869__A2 _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09664_ _00118_ io_in[4] u_cpu.rf_ram.memory\[45\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06876_ _02959_ _03002_ _03005_ _00353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05424__S0 _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05827_ u_cpu.cpu.bufreg2.i_cnt_done _02311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08615_ u_arbiter.i_wb_cpu_dbus_adr\[28\] u_arbiter.i_wb_cpu_dbus_adr\[27\] _04115_
+ _04130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09595_ _00049_ io_in[4] u_cpu.rf_ram.memory\[81\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06541__A2 _02812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08818__A1 _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05758_ _02236_ _02238_ _02240_ _02242_ _01425_ _02243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_08546_ u_cpu.rf_ram.memory\[31\]\[0\] _04094_ _04095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08818__B2 _04024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08477_ _03747_ _03988_ _03801_ _04040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09737__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09491__A1 _04468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08294__A2 _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05689_ _01594_ _02174_ _01626_ _02175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08483__B _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05727__S1 _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07428_ u_cpu.rf_ram.memory\[132\]\[7\] _03305_ _03313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_u_scanchain_local.scan_flop\[41\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10714__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07359_ _03274_ _03275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08046__A2 _03654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06057__A1 _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09887__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10370_ _00803_ io_in[4] u_cpu.rf_ram.memory\[11\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09029_ _02810_ _04197_ _04378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[56\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10864__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09546__A2 _04674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05032__A2 _01457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07309__A1 _03161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06780__A2 _02944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06532__A2 _02801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10244__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08809__A1 _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10706_ _01135_ io_in[4] u_cpu.rf_ram.memory\[104\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10394__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10637_ _01066_ io_in[4] u_cpu.rf_ram.memory\[94\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09234__A1 _04484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10568_ _00998_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08613__S _04115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07796__A1 _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06599__A2 _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10499_ _00932_ io_in[4] u_cpu.rf_ram.memory\[32\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09537__A2 _04664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05271__A2 _01761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07548__A1 _03343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_04991_ u_arbiter.i_wb_cpu_dbus_adr\[18\] _01442_ _01497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06771__A2 _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06730_ _02750_ _02914_ _02920_ _00292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06661_ u_cpu.rf_ram.memory\[76\]\[7\] _02874_ _02882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06523__A2 _02801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05612_ _01422_ _02089_ _02098_ _02099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_08400_ _01436_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[9\] _03972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__07899__S _03586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09380_ _02311_ _02344_ _01386_ _04581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_36_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06592_ _02843_ _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08331_ _03907_ _03909_ _03911_ _03876_ _03912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_33_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10737__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05543_ _01539_ _02021_ _02030_ _02031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__08276__A2 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05720__B _01402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08262_ _03847_ _03850_ _03852_ _03853_ _03854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_05474_ u_cpu.rf_ram.memory\[0\]\[4\] u_cpu.rf_ram.memory\[1\]\[4\] u_cpu.rf_ram.memory\[2\]\[4\]
+ u_cpu.rf_ram.memory\[3\]\[4\] _01556_ _01557_ _01962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07213_ u_cpu.rf_ram.memory\[71\]\[7\] _03186_ _03194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08193_ _03752_ _03771_ _03783_ _03792_ _03793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_20_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06039__A1 _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07144_ _03152_ _00474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10887__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07075_ _03114_ _00443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09528__A2 _04664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06026_ u_cpu.rf_ram.memory\[82\]\[0\] _02477_ _02483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07139__S _03148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10117__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07977_ u_cpu.rf_ram.memory\[116\]\[3\] _03626_ _03630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06762__A2 _02934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10267__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09716_ _00170_ io_in[4] u_cpu.rf_ram.memory\[50\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_101_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06928_ u_cpu.rf_ram.memory\[58\]\[2\] _03031_ _03034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09647_ _00101_ io_in[4] u_cpu.rf_ram.memory\[42\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06859_ u_cpu.rf_ram.memory\[61\]\[3\] _02992_ _02996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06514__A2 _02791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09578_ _00032_ io_in[4] u_cpu.rf_ram.memory\[82\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08529_ _03539_ _04084_ _04085_ _00927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08267__A2 _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09464__A1 _04478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06278__A1 _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09216__A1 _04484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10422_ _00855_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07078__I0 _02596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07778__A1 _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10353_ _00786_ io_in[4] u_cpu.rf_ram.memory\[121\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07049__S _03100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06450__A1 _02754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09519__A2 _04654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10284_ _00717_ io_in[4] u_cpu.rf_ram.memory\[91\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08727__B1 _04175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07950__A1 _03555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06753__A2 _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09902__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05805__B _01648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06505__A2 _02791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09207__A1 _04478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05190_ u_cpu.rf_ram.memory\[136\]\[0\] u_cpu.rf_ram.memory\[137\]\[0\] u_cpu.rf_ram.memory\[138\]\[0\]
+ u_cpu.rf_ram.memory\[139\]\[0\] _01680_ _01681_ _01682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_127_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08430__A2 u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06441__A1 _02748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08718__B1 _04175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06992__A2 _03061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07900_ _03587_ _00796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08880_ _02516_ _04296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_123_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08194__A1 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07831_ u_cpu.rf_ram.memory\[120\]\[3\] _03541_ _03548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09582__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06744__A2 _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07762_ _03357_ _03500_ _03507_ _00738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_04974_ u_cpu.cpu.ctrl.o_ibus_adr\[14\] _01481_ _01442_ _01484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09501_ _04480_ _04644_ _04650_ _01334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06713_ u_cpu.rf_ram.memory\[68\]\[6\] _02904_ _02911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07693_ _03464_ _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_65_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06644_ _02754_ _02864_ _02872_ _00254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_64_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09432_ _04482_ _04605_ _04612_ _01303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09363_ _04567_ _04568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06575_ u_cpu.rf_ram.memory\[129\]\[0\] _02834_ _02835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05180__A1 _01553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09446__A1 _04478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05526_ _01398_ _02013_ _02014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08314_ _03890_ _03891_ _03894_ _03895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09294_ u_cpu.rf_ram.memory\[86\]\[2\] _04526_ _04529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08245_ _03773_ _03767_ _03801_ _03838_ _03811_ _03839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_05457_ u_cpu.rf_ram.memory\[136\]\[3\] u_cpu.rf_ram.memory\[137\]\[3\] u_cpu.rf_ram.memory\[138\]\[3\]
+ u_cpu.rf_ram.memory\[139\]\[3\] _01680_ _01681_ _01946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_20_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06680__A1 _02754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08176_ _03775_ _03776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05388_ _01870_ _01872_ _01874_ _01876_ _01568_ _01877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_118_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07127_ _02961_ _03139_ _03143_ _00466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08421__A2 _03985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06432__A1 _02742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07058_ _03105_ _00435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_79_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06009_ _01543_ _02465_ _02466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06983__A2 _03061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09925__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08185__A1 _02765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07932__A1 _03555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06735__A2 _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10902__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05094__S1 _01580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05625__B _01565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10971_ _10971_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_44_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07160__A2 _03159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05171__A1 _01609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[60\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08660__A2 _04155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08163__S _01435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10405_ _00838_ io_in[4] u_cpu.rf_ram.memory\[33\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10432__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07471__I0 _02584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10336_ _00769_ io_in[4] u_cpu.rf_ram.memory\[120\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06974__A2 _03051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10267_ _00700_ io_in[4] u_cpu.rf_ram.memory\[36\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04985__A1 _01443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05609__S0 _01623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10198_ _00644_ io_in[4] u_cpu.rf_ram.memory\[127\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10582__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06726__A2 _02914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08971__I0 u_arbiter.i_wb_cpu_rdt\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08479__A2 _03818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09428__A1 _04478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06360_ _02497_ _02697_ _02701_ _00141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08100__A1 u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05311_ _01589_ _01800_ _01801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06291_ _02521_ _02624_ _02660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08651__A2 _04145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08030_ _03667_ _00846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_05242_ u_cpu.rf_ram.memory\[108\]\[1\] u_cpu.rf_ram.memory\[109\]\[1\] u_cpu.rf_ram.memory\[110\]\[1\]
+ u_cpu.rf_ram.memory\[111\]\[1\] _01619_ _01620_ _01733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06662__A1 _02754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05173_ _01553_ _01664_ _01654_ _01665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09948__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06414__A1 _02492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09981_ _00435_ io_in[4] u_cpu.rf_ram.memory\[9\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05768__A3 _02252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06965__A2 _03051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10925__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08932_ u_cpu.rf_ram.memory\[28\]\[3\] _04322_ _04326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08167__A1 _02765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08863_ u_cpu.rf_ram.memory\[94\]\[1\] _04282_ _04285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06717__A2 _02682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07814_ _03355_ _03530_ _03536_ _00761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08794_ u_cpu.rf_ram.memory\[93\]\[5\] _04227_ _04233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07390__A2 _03285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05164__C _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04957_ _01470_ _01464_ _01471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07745_ u_cpu.cpu.state.init_done _03458_ _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04888_ u_cpu.cpu.immdec.imm24_20\[1\] _01387_ _01413_ _01414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07676_ _01428_ _03453_ _03454_ _00704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_80_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10305__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09415_ u_cpu.rf_ram.memory\[27\]\[7\] _04595_ _04603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06627_ _02626_ _02638_ _02863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08890__A2 _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05180__B _01565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09346_ u_cpu.rf_ram.memory\[88\]\[1\] _04556_ _04558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06558_ u_cpu.rf_ram.memory\[119\]\[1\] _02823_ _02825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05509_ _01594_ _01996_ _01416_ _01997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09277_ _04474_ _04516_ _04519_ _01241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06489_ u_cpu.rf_ram_if.rcnt\[0\] _02784_ _00187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_32_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08642__A2 _04145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10455__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08228_ _01374_ _02768_ _03824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_5_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08159_ _02765_ u_arbiter.i_wb_cpu_rdt\[5\] _03758_ _03759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_134_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06405__A1 _02517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10121_ _00567_ io_in[4] u_cpu.rf_ram.memory\[135\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06956__A2 _03041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08158__A1 _01436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10052_ _00498_ io_in[4] u_cpu.rf_ram.memory\[71\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06708__A2 _02904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08953__I0 u_arbiter.i_wb_cpu_rdt\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_u_scanchain_local.scan_flop\[8\]_SI u_arbiter.i_wb_cpu_dbus_dat\[2\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07381__A2 _03285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05392__A1 _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10954_ u_cpu.cpu.o_wdata1 io_in[4] u_cpu.rf_ram_if.wdata1_r\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08330__A1 _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07133__A2 _03139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08881__A2 _04282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10885_ _01314_ io_in[4] u_cpu.rf_ram.memory\[24\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06892__A1 _02957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08094__B1 _03654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[65\] u_scanchain_local.module_data_in\[64\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[27\] u_scanchain_local.clk u_scanchain_local.module_data_in\[65\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_89_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06644__A1 _02754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05447__A2 _01935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10948__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08397__A1 _03762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06947__A2 _03041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10319_ _00752_ io_in[4] u_cpu.rf_ram.memory\[34\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05860_ u_cpu.cpu.decode.op21 _02343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09361__A3 _02338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07372__A2 _03275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10328__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05791_ u_cpu.rf_ram.memory\[88\]\[7\] u_cpu.rf_ram.memory\[89\]\[7\] u_cpu.rf_ram.memory\[90\]\[7\]
+ u_cpu.rf_ram.memory\[91\]\[7\] _01646_ _01603_ _02276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__05383__A1 _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07530_ _03343_ _03372_ _03373_ _00639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_93_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09620__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08321__A1 _03742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07124__A2 _03139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07461_ _03169_ _03325_ _03331_ _00612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05135__A1 _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08872__A2 _04282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06412_ _02487_ _02729_ _02731_ _00163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09200_ u_cpu.rf_ram.memory\[84\]\[2\] _04470_ _04475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10478__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07392_ u_cpu.rf_ram.memory\[134\]\[7\] _03285_ _03293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09131_ u_cpu.rf_ram.memory\[107\]\[5\] _04429_ _04435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06343_ _02502_ _02686_ _02691_ _00134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08624__A2 _02448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09770__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09062_ _04294_ _04389_ _04396_ _01149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06274_ _02650_ _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08013_ _03652_ _03653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05225_ _01594_ _01715_ _01564_ _01716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08388__A1 _03756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05156_ _01416_ _01648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_143_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06938__A2 _03031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09964_ _00418_ io_in[4] u_cpu.rf_ram.memory\[53\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05087_ _01547_ _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07147__S _03148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08915_ u_cpu.rf_ram.memory\[96\]\[6\] _04309_ _04316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09895_ _00349_ io_in[4] u_cpu.rf_ram.memory\[61\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08846_ _03545_ _04271_ _04274_ _01055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07363__A2 _03275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05213__I2 u_cpu.rf_ram.memory\[22\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05374__A1 _01399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08777_ _04223_ _01037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05989_ _02450_ _02451_ _02449_ _00023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_84_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07728_ _02432_ _02434_ _03484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08312__A1 _03831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07115__A2 _03129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05126__A1 _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07659_ u_cpu.rf_ram.memory\[36\]\[2\] _03442_ _03445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06174__I0 _02587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08863__A2 _04282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06874__A1 _02957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10670_ _01099_ io_in[4] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09329_ _04472_ _04546_ _04548_ _01264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06626__A1 _02754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08379__A1 _03797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06025__I _02481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09040__A2 _04379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06929__A2 _03031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07057__S _03100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05601__A2 _02087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10104_ _00550_ io_in[4] u_cpu.rf_ram.memory\[137\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11084_ _11084_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_89_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10035_ _00481_ io_in[4] u_cpu.rf_ram.memory\[72\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09643__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07354__A2 _03265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08551__A1 _03545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05365__A1 _01636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10620__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07106__A2 _03129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10937_ u_cpu.rf_ram_if.wdata0_r\[4\] io_in[4] u_cpu.rf_ram_if.wdata0_r\[3\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08854__A2 _04271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09793__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10868_ _01297_ io_in[4] u_cpu.rf_ram.memory\[26\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08067__B1 _03678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10770__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10799_ _01228_ io_in[4] u_cpu.rf_ram.memory\[10\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06093__A2 _02530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07290__A1 u_cpu.rf_ram.memory\[39\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10000__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05010_ u_cpu.cpu.ctrl.o_ibus_adr\[23\] _01509_ _01511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_126_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09031__A2 _04379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07593__A2 _03402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10150__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06961_ _02953_ _03051_ _03052_ _00391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08700_ u_cpu.cpu.ctrl.o_ibus_adr\[20\] _04173_ _04175_ u_cpu.cpu.ctrl.o_ibus_adr\[21\]
+ _04180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05912_ _02311_ _02315_ _02316_ _02393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_09680_ _00134_ io_in[4] u_cpu.rf_ram.memory\[51\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06892_ _02957_ _03012_ _03014_ _00360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07345__A2 _03265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08631_ _02361_ _04139_ _04140_ _00974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05356__A1 _01553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05843_ _02309_ u_cpu.cpu.alu.add_cy_r _02327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08562_ u_cpu.cpu.alu.cmp_r _02433_ _04103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09098__A2 _04409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05774_ u_cpu.rf_ram.memory\[100\]\[7\] u_cpu.rf_ram.memory\[101\]\[7\] u_cpu.rf_ram.memory\[102\]\[7\]
+ u_cpu.rf_ram.memory\[103\]\[7\] _01577_ _01549_ _02259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_82_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07513_ u_cpu.rf_ram.memory\[128\]\[1\] _03362_ _03364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05108__A1 _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08493_ _03973_ _04028_ _04054_ _03851_ _04055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_126_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08845__A2 _04271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06856__A1 _02957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07444_ u_cpu.rf_ram.memory\[131\]\[6\] _03315_ _03322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08058__B1 _03678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07375_ _03173_ _03275_ _03283_ _00574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09114_ _04292_ _04419_ _04425_ _01172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06608__A1 _02754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06326_ _02512_ _02673_ _02680_ _00128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09270__A2 _04197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09045_ u_cpu.rf_ram.memory\[104\]\[7\] _04379_ _04387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06257_ u_cpu.rf_ram.memory\[42\]\[0\] _02641_ _02642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06084__A2 _02530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07281__A1 _03169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05208_ u_cpu.rf_ram.memory\[4\]\[1\] u_cpu.rf_ram.memory\[5\]\[1\] u_cpu.rf_ram.memory\[6\]\[1\]
+ u_cpu.rf_ram.memory\[7\]\[1\] _01546_ _01550_ _01699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_11_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05831__A2 _02312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06188_ u_cpu.rf_ram_if.wdata1_r\[7\] u_cpu.cpu.o_wdata0 _02460_ _02598_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09022__A2 _04369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07033__A1 _02953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05139_ _01539_ _01569_ _01588_ _01630_ _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_143_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09666__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07584__A2 _03402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09947_ _00401_ io_in[4] u_cpu.rf_ram.memory\[55\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05595__A1 _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10643__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09878_ _00332_ io_in[4] u_cpu.rf_ram.memory\[63\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08533__A1 _03545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07336__A2 _03255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08829_ u_cpu.cpu.immdec.imm11_7\[3\] _04236_ _04262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05347__B2 _01836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09089__A2 _04409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10793__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08836__A2 _03741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10722_ _01151_ io_in[4] u_cpu.rf_ram.memory\[79\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10653_ _01082_ io_in[4] u_cpu.rf_ram.memory\[96\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10023__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10584_ _01014_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09261__A2 _04506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09013__A2 _04369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10173__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05808__B _01402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[28\] u_arbiter.i_wb_cpu_rdt\[25\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[22\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__07575__A2 _03392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05586__A1 _01397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11067_ _11067_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_27_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07327__A2 _03255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10018_ _00464_ io_in[4] u_cpu.rf_ram.memory\[140\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05433__S1 _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08827__A2 _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06838__A1 _02957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07886__I0 _02584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05490_ u_cpu.rf_ram.memory\[60\]\[4\] u_cpu.rf_ram.memory\[61\]\[4\] u_cpu.rf_ram.memory\[62\]\[4\]
+ u_cpu.rf_ram.memory\[63\]\[4\] _01598_ _01573_ _01978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08346__S _01436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05197__S0 _01687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07160_ _03161_ _03159_ _03162_ _00480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09252__A2 _02524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06111_ u_cpu.rf_ram.memory\[81\]\[5\] _02541_ _02547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10516__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07091_ _02961_ _03119_ _03123_ _00450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09689__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06042_ _02495_ _02496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09004__A2 _04359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07015__A1 _02953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10666__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07566__A2 _03392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09801_ _00255_ io_in[4] u_cpu.rf_ram.memory\[76\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05577__A1 _01540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07993_ u_cpu.rf_ram.memory\[33\]\[2\] _03636_ _03639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09732_ _00186_ io_in[4] u_cpu.rf_ram_if.rreq_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06944_ u_cpu.rf_ram.memory\[57\]\[1\] _03041_ _03043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08515__A1 _01374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07318__A2 _03245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09663_ _00117_ io_in[4] u_cpu.rf_ram.memory\[45\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05329__A1 _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06875_ u_cpu.rf_ram.memory\[60\]\[2\] _03002_ _03005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05453__B _01417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08614_ _04129_ _00968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05424__S1 _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05826_ _02309_ u_cpu.cpu.alu.add_cy_r _02310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09594_ _00048_ io_in[4] u_cpu.rf_ram.memory\[81\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08545_ _04093_ _04094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_54_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05757_ _01601_ _02241_ _01605_ _02242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_23_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10046__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08476_ _03788_ _03776_ _03851_ _03896_ _04039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_05688_ u_cpu.rf_ram.memory\[96\]\[6\] u_cpu.rf_ram.memory\[97\]\[6\] u_cpu.rf_ram.memory\[98\]\[6\]
+ u_cpu.rf_ram.memory\[99\]\[6\] _01602_ _01579_ _02174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_50_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09491__A2 _04644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07427_ _03171_ _03305_ _03312_ _00597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07358_ _02602_ _02832_ _03274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10196__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06309_ _02517_ _02662_ _02670_ _00121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06057__A2 _02507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07289_ _03157_ _03235_ _03236_ _00535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09028_ _04296_ _04369_ _04377_ _01134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05360__S0 _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07557__A2 _03382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[17\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05347__C _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05568__A1 _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05112__S0 _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08506__A1 _04016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07309__A2 _03245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05179__S0 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07070__S _03109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10539__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06296__A2 _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10705_ _01134_ io_in[4] u_cpu.rf_ram.memory\[103\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07493__A1 _03349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10636_ _01065_ io_in[4] u_cpu.rf_ram.memory\[94\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09831__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[31\]_D u_arbiter.i_wb_cpu_rdt\[28\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09234__A2 _04487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10567_ _00997_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10689__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07796__A2 _03520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08993__A1 _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10498_ _00931_ io_in[4] u_cpu.rf_ram.memory\[32\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05351__S0 _01646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09981__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07548__A2 _03382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08745__A1 _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05559__A1 _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05103__S0 _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06220__A2 _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04990_ u_cpu.cpu.ctrl.o_ibus_adr\[17\] _01491_ u_cpu.cpu.ctrl.o_ibus_adr\[18\] _01496_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_77_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09170__A1 _04294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10069__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05273__B _01565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06660_ _02752_ _02874_ _02881_ _00261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07720__A2 _03475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05611_ _02091_ _02093_ _02095_ _02097_ _01607_ _02098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05731__A1 _01406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06591_ _02706_ _02832_ _02843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08330_ _03780_ _03910_ _03911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05542_ _02023_ _02025_ _02027_ _02029_ _01568_ _02030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_71_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06287__A2 _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08261_ _02768_ _03774_ _03853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05473_ _01554_ _01960_ _01961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07484__A1 _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07212_ _03171_ _03186_ _03193_ _00501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08192_ _03786_ _03790_ _03791_ _03792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09225__A2 _04487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06039__A2 _02492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07236__A1 _03157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07143_ _02587_ u_cpu.rf_ram.memory\[13\]\[3\] _03148_ _03152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07787__A2 _03520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08984__A1 _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07074_ _02590_ u_cpu.rf_ram.memory\[15\]\[4\] _03109_ _03114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_126_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06025_ _02481_ _02482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07539__A2 _03372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07976_ _03545_ _03626_ _03629_ _00830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09715_ _00169_ io_in[4] u_cpu.rf_ram.memory\[47\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06927_ _02957_ _03031_ _03033_ _00376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09704__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09646_ _00100_ io_in[4] u_cpu.rf_ram.memory\[42\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06858_ _02959_ _02992_ _02995_ _00345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05809_ u_cpu.rf_ram.memory\[136\]\[7\] u_cpu.rf_ram.memory\[137\]\[7\] u_cpu.rf_ram.memory\[138\]\[7\]
+ u_cpu.rf_ram.memory\[139\]\[7\] _01687_ _01688_ _02294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09577_ _00031_ io_in[4] u_cpu.rf_ram.memory\[82\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05722__A1 _01399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06789_ _02481_ _02953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08528_ u_cpu.rf_ram.memory\[32\]\[0\] _04084_ _04085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09854__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09464__A2 _04625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06278__A2 _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08672__B1 _04157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08459_ _03845_ _04022_ _04023_ _00919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__05630__C _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10831__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[13\]_D u_arbiter.i_wb_cpu_rdt\[10\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09216__A2 _04470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10421_ _00854_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07778__A2 _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08975__A1 _02524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10352_ _00785_ io_in[4] u_cpu.rf_ram.memory\[121\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06450__A2 _02740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10283_ _00716_ io_in[4] u_cpu.rf_ram.memory\[91\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08727__B2 _04195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05077__C _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10211__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05261__I0 u_cpu.rf_ram.memory\[92\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07950__A2 _03606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05961__A1 _01403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09152__A1 _04294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07702__A2 _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10361__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05713__A1 _01553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09455__A2 _04625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06269__A2 _02641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07466__A1 _02577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09207__A2 _04470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07218__A1 _03157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10619_ _01048_ io_in[4] u_cpu.cpu.immdec.imm11_7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07769__A2 _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05268__B _01654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06441__A2 _02740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09727__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08194__A2 _03793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07830_ _02496_ _03547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[40\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07941__A2 _03606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07761_ u_cpu.rf_ram.memory\[92\]\[6\] _03500_ _03507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_04973_ u_arbiter.i_wb_cpu_dbus_adr\[14\] _01443_ _01483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10704__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09500_ u_cpu.rf_ram.memory\[98\]\[5\] _04644_ _04650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06712_ _02750_ _02904_ _02910_ _00284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07692_ _02475_ _02706_ _03464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09877__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09431_ u_cpu.rf_ram.memory\[26\]\[6\] _04605_ _04612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06643_ u_cpu.rf_ram.memory\[74\]\[7\] _02864_ _02872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05704__A1 _01645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[55\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09362_ _04565_ _04566_ _04567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__10854__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06574_ _02833_ _02834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09446__A2 _04615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08313_ _03893_ _03894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05525_ u_cpu.rf_ram.memory\[92\]\[4\] u_cpu.rf_ram.memory\[93\]\[4\] u_cpu.rf_ram.memory\[94\]\[4\]
+ u_cpu.rf_ram.memory\[95\]\[4\] _01610_ _01611_ _02013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_61_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07457__A1 _03165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09293_ _04472_ _04526_ _04528_ _01248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08244_ _03761_ _03790_ _03835_ _03837_ _03838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_05456_ _01925_ _01944_ _01402_ _01945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06680__A2 _02884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08175_ u_arbiter.i_wb_cpu_rdt\[14\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[14\]
+ _01435_ _03775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05387_ _01562_ _01875_ _01565_ _01876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_10_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07126_ u_cpu.rf_ram.memory\[140\]\[3\] _03139_ _03143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07057_ _02590_ u_cpu.rf_ram.memory\[9\]\[4\] _03100_ _03105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06432__A2 _02740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10234__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06008_ u_cpu.rf_ram_if.rcnt\[1\] u_cpu.rf_ram_if.rcnt\[0\] u_cpu.rf_ram_if.rcnt\[2\]
+ _02465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_115_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08185__A2 u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07932__A2 _03596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10384__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07959_ u_cpu.rf_ram.memory\[115\]\[3\] _03616_ _03620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05943__A1 _02320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09134__A1 _04294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10970_ _10970_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_16_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09629_ _00083_ io_in[4] u_cpu.rf_ram.memory\[80\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09437__A2 _04615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07448__A1 _02469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07999__A2 _03636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06120__A1 _02482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06671__A2 _02884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06472__B _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10404_ _00837_ io_in[4] u_cpu.rf_ram.memory\[33\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10335_ _00768_ io_in[4] u_cpu.rf_ram.memory\[120\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06423__A2 _02729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07620__A1 _03343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10266_ _00699_ io_in[4] u_cpu.rf_ram.memory\[36\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08399__B _03906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10727__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[10\] u_arbiter.i_wb_cpu_rdt\[7\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[4\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__05609__S1 _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05816__B _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10197_ _00643_ io_in[4] u_cpu.rf_ram.memory\[127\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07923__A2 _03596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05934__A1 _02320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08619__S _02372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10877__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07687__A1 _01429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05793__S0 _01590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09428__A2 _04605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10107__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07439__A1 _03165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08100__A2 _03654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05310_ u_cpu.rf_ram.memory\[52\]\[2\] u_cpu.rf_ram.memory\[53\]\[2\] u_cpu.rf_ram.memory\[54\]\[2\]
+ u_cpu.rf_ram.memory\[55\]\[2\] _01590_ _01591_ _01800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_06290_ _02517_ _02651_ _02659_ _00113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05545__S0 _01680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05241_ _01539_ _01703_ _01712_ _01731_ _01732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__06662__A2 _02874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10257__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08939__A1 _04294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05172_ u_cpu.rf_ram.memory\[84\]\[0\] u_cpu.rf_ram.memory\[85\]\[0\] u_cpu.rf_ram.memory\[86\]\[0\]
+ u_cpu.rf_ram.memory\[87\]\[0\] _01555_ _01652_ _01664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_122_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06414__A2 _02729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09980_ _00434_ io_in[4] u_cpu.rf_ram.memory\[9\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08931_ _04286_ _04322_ _04325_ _01089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08167__A2 u_arbiter.i_wb_cpu_rdt\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09364__A1 u_cpu.cpu.genblk3.csr.o_new_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08862_ _02486_ _04284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07813_ u_cpu.rf_ram.memory\[117\]\[5\] _03530_ _03536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08793_ _03549_ _04227_ _04232_ _01044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05445__C _01426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09116__A1 _04294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07744_ _03497_ _00730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_04956_ u_cpu.cpu.ctrl.o_ibus_adr\[9\] _01470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_26_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07678__A1 u_cpu.cpu.mem_bytecnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07675_ u_cpu.cpu.state.o_cnt\[2\] u_cpu.cpu.state.o_cnt_r\[3\] _03454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_04887_ _01411_ _01412_ u_cpu.rf_ram_if.rtrig0 _01377_ _01413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_77_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09414_ _04482_ _04595_ _04602_ _01295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06626_ _02754_ _02854_ _02862_ _00246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09419__A2 _04605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09345_ _04468_ _04556_ _04557_ _01271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06557_ _02738_ _02823_ _02824_ _00215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08627__B1 _04137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05508_ u_cpu.rf_ram.memory\[104\]\[4\] u_cpu.rf_ram.memory\[105\]\[4\] u_cpu.rf_ram.memory\[106\]\[4\]
+ u_cpu.rf_ram.memory\[107\]\[4\] _01615_ _01616_ _01996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_138_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09276_ u_cpu.rf_ram.memory\[110\]\[2\] _04516_ _04519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06102__A1 _02482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05536__S0 _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06488_ _02769_ _02783_ _02784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08227_ _03823_ _00887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_138_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05439_ u_cpu.rf_ram.memory\[88\]\[3\] u_cpu.rf_ram.memory\[89\]\[3\] u_cpu.rf_ram.memory\[90\]\[3\]
+ u_cpu.rf_ram.memory\[91\]\[3\] _01646_ _01603_ _01928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07850__A1 _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06653__A2 _02874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08158_ _01436_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[5\] _03758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_134_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07109_ _02961_ _03129_ _03133_ _00458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07602__A1 _03343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06405__A2 _02718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08089_ u_arbiter.i_wb_cpu_rdt\[20\] _03669_ _03654_ u_arbiter.i_wb_cpu_dbus_dat\[20\]
+ _03709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_122_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10120_ _00566_ io_in[4] u_cpu.rf_ram.memory\[136\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04967__A2 _01457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09355__A1 _04480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05636__B _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10051_ _00497_ io_in[4] u_cpu.rf_ram.memory\[71\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05916__A1 u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05392__A2 _01880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10953_ u_cpu.rf_ram_if.wdata1_r\[7\] io_in[4] u_cpu.rf_ram_if.wdata1_r\[6\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06341__A1 _02497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10884_ _01313_ io_in[4] u_cpu.rf_ram.memory\[24\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06892__A2 _03012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08094__A1 u_arbiter.i_wb_cpu_rdt\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05527__S0 _01646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07141__I0 _02584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09572__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07841__A1 _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06644__A2 _02864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[58\] u_scanchain_local.module_data_in\[57\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[20\] u_scanchain_local.clk u_scanchain_local.module_data_in\[58\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_106_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10318_ _00751_ io_in[4] u_cpu.rf_ram.memory\[34\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10249_ _00682_ io_in[4] u_cpu.rf_ram.memory\[38\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05907__A1 _01369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05790_ _01398_ _02274_ _02275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05383__A2 _01871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06580__A1 _02744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07460_ u_cpu.rf_ram.memory\[130\]\[5\] _03325_ _03331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06332__A1 _02682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06411_ u_cpu.rf_ram.memory\[47\]\[1\] _02729_ _02731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06883__A2 _03002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07391_ _03171_ _03285_ _03292_ _00581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09915__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09130_ _04290_ _04429_ _04434_ _01179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06342_ u_cpu.rf_ram.memory\[51\]\[4\] _02686_ _02691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09061_ u_cpu.rf_ram.memory\[99\]\[6\] _04389_ _04396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07832__A1 _03547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06273_ _02625_ _02639_ _02650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06635__A2 _02864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08012_ u_arbiter.i_wb_cpu_ack _01442_ _03652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_135_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05224_ u_cpu.rf_ram.memory\[48\]\[1\] u_cpu.rf_ram.memory\[49\]\[1\] u_cpu.rf_ram.memory\[50\]\[1\]
+ u_cpu.rf_ram.memory\[51\]\[1\] _01544_ _01548_ _01715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_128_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08388__A2 _03810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05155_ u_cpu.rf_ram.memory\[120\]\[0\] u_cpu.rf_ram.memory\[121\]\[0\] u_cpu.rf_ram.memory\[122\]\[0\]
+ u_cpu.rf_ram.memory\[123\]\[0\] _01646_ _01603_ _01647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_144_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06399__A1 _02502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09963_ _00417_ io_in[4] u_cpu.rf_ram.memory\[53\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05086_ _01577_ _01578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09337__A1 _04480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08914_ _04292_ _04309_ _04315_ _01082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05456__B _01402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09894_ _00348_ io_in[4] u_cpu.rf_ram.memory\[61\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[50\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08845_ u_cpu.rf_ram.memory\[97\]\[2\] _04271_ _04274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08560__A2 _04094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08776_ _02593_ u_cpu.rf_ram.memory\[2\]\[5\] _04217_ _04223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06571__A1 _02754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05970__I _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05988_ _02379_ _02380_ _02451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07727_ _03359_ _03475_ _03483_ _00726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04939_ _01442_ _01457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10422__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07658_ _03347_ _03442_ _03444_ _00696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05126__A2 _01617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06609_ _02626_ _02660_ _02853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09595__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06874__A2 _03002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07589_ u_cpu.rf_ram.memory\[124\]\[3\] _03402_ _03406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04885__A1 _01410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09328_ u_cpu.rf_ram.memory\[87\]\[1\] _04546_ _04548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10572__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07823__A1 _03539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06626__A2 _02854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09259_ _04474_ _04506_ _04509_ _01233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10103_ _00549_ io_in[4] u_cpu.rf_ram.memory\[137\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11083_ _11083_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_49_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08000__A1 _03551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10034_ _00480_ io_in[4] u_cpu.rf_ram.memory\[72\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[3\] u_arbiter.i_wb_cpu_rdt\[0\] io_in[3] u_arbiter.i_wb_cpu_dbus_sel\[1\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__08551__A2 _04094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06562__A1 u_cpu.rf_ram.memory\[119\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09938__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08303__A2 _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10936_ u_cpu.rf_ram_if.wdata0_r\[3\] io_in[4] u_cpu.rf_ram_if.wdata0_r\[2\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06314__A1 _02482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10915__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06865__A2 _02992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10867_ _01296_ io_in[4] u_cpu.rf_ram.memory\[27\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08067__A1 u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10798_ _01227_ io_in[4] u_cpu.rf_ram.memory\[10\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07814__A1 _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06617__A2 _02854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07290__A2 _03235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09567__A1 _01429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07042__A2 _03091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09319__A1 _04480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08790__A2 _04227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06960_ u_cpu.rf_ram.memory\[56\]\[0\] _03051_ _03052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05911_ u_cpu.cpu.immdec.imm31 _02317_ _02392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_67_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06891_ u_cpu.rf_ram.memory\[19\]\[1\] _03012_ _03014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08542__A2 _04084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08630_ u_cpu.cpu.bufreg.lsb\[1\] _04139_ _04140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10445__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05842_ _02308_ _02325_ _02326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__05356__A2 _01845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08561_ _03555_ _04094_ _04102_ _00942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05773_ _01594_ _02257_ _01416_ _02258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07512_ _03343_ _03362_ _03363_ _00631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06305__A1 _02507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08492_ _04024_ _04053_ _04054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05108__A2 _01599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10595__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07443_ _03169_ _03315_ _03321_ _00604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06856__A2 _02992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04867__A1 u_cpu.cpu.genblk3.csr.o_new_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08058__A1 u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07374_ u_cpu.rf_ram.memory\[135\]\[7\] _03275_ _03283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09113_ u_cpu.rf_ram.memory\[106\]\[5\] _04419_ _04425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06325_ u_cpu.rf_ram.memory\[44\]\[6\] _02673_ _02680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06608__A2 _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09044_ _04294_ _04379_ _04386_ _01141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06256_ _02640_ _02641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07281__A2 _03225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05207_ _01554_ _01697_ _01417_ _01698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_85_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08605__I0 u_arbiter.i_wb_cpu_dbus_adr\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06187_ _02597_ _00072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08230__A1 _03754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07033__A2 _03091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05138_ _01422_ _01608_ _01629_ _01630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_89_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05069_ _01554_ _01560_ _01561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09946_ _00400_ io_in[4] u_cpu.rf_ram.memory\[55\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05595__A2 _02081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06792__A1 u_cpu.rf_ram.memory\[29\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09877_ _00331_ io_in[4] u_cpu.rf_ram.memory\[63\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08533__A2 _04084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08828_ _03801_ _03900_ _04260_ _04261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06544__A1 _02746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08759_ _02593_ u_cpu.rf_ram.memory\[3\]\[5\] _04208_ _04214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_57_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10938__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10721_ _01150_ io_in[4] u_cpu.rf_ram.memory\[99\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06847__A2 _02982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10652_ _01081_ io_in[4] u_cpu.rf_ram.memory\[96\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10583_ _01013_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07272__A2 _03225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10318__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09549__A1 _04474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07068__S _03109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08221__A1 _03769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07024__A2 _03081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09610__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10468__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05586__A2 _02072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11066_ _11066_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_114_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09760__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10017_ _00463_ io_in[4] u_cpu.rf_ram.memory\[140\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06535__A1 _02639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08288__A1 _02337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05115__I _01425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10919_ _01348_ io_in[4] u_cpu.rf_ram.memory\[89\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06838__A2 _02982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05197__S1 _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06110_ _02502_ _02541_ _02546_ _00046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08460__A1 _03973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07090_ u_cpu.rf_ram.memory\[142\]\[3\] _03119_ _03123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06041_ _02460_ u_cpu.rf_ram_if.wdata0_r\[3\] _02494_ _02495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07015__A2 _03081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05718__C _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09800_ _00254_ io_in[4] u_cpu.rf_ram.memory\[74\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07992_ _03543_ _03636_ _03638_ _00837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05577__A2 _02063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06774__A1 _02738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09731_ _00185_ io_in[4] u_cpu.rf_ram.memory\[4\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06943_ _02953_ _03041_ _03042_ _00383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09662_ _00116_ io_in[4] u_cpu.rf_ram.memory\[45\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06874_ _02957_ _03002_ _03004_ _00352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05329__A2 _01790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08613_ u_arbiter.i_wb_cpu_dbus_adr\[27\] u_arbiter.i_wb_cpu_dbus_adr\[26\] _04115_
+ _04129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05825_ u_cpu.cpu.alu.i_rs1 _02309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09593_ _00047_ io_in[4] u_cpu.rf_ram.memory\[81\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08544_ _02528_ _02727_ _04093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05756_ u_cpu.rf_ram.memory\[56\]\[7\] u_cpu.rf_ram.memory\[57\]\[7\] u_cpu.rf_ram.memory\[58\]\[7\]
+ u_cpu.rf_ram.memory\[59\]\[7\] _01602_ _01579_ _02241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_70_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08475_ _03779_ _04037_ _04038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06829__A2 _02972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05687_ _01636_ _02172_ _02173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07426_ u_cpu.rf_ram.memory\[132\]\[6\] _03305_ _03312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07357_ _03173_ _03265_ _03273_ _00566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06308_ u_cpu.rf_ram.memory\[45\]\[7\] _02662_ _02670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09633__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07288_ u_cpu.rf_ram.memory\[39\]\[0\] _03235_ _03236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09027_ u_cpu.rf_ram.memory\[103\]\[7\] _04369_ _04377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06239_ _02487_ _02628_ _02630_ _00091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05360__S1 _01652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10610__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07006__A2 _03071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05017__A1 _01445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09783__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05568__A2 _02054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05112__S1 _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09929_ _00383_ io_in[4] u_cpu.rf_ram.memory\[57\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10760__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07190__A1 _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05740__A2 _02220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05179__S1 _01549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10704_ _01133_ io_in[4] u_cpu.rf_ram.memory\[103\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07493__A2 _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10140__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10635_ _01064_ io_in[4] u_cpu.rf_ram.memory\[94\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08442__A1 _02433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10566_ _00996_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07245__A2 _03206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05256__A1 _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08993__A2 _04197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[40\] u_scanchain_local.module_data_in\[39\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[2\] u_scanchain_local.clk u_scanchain_local.module_data_in\[40\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
X_10497_ _00930_ io_in[4] u_cpu.rf_ram.memory\[32\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10290__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05351__S1 _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09242__I0 _02587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08745__A2 _04199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05103__S1 _01548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06756__A1 _02738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11049_ _11049_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_37_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09170__A2 _04449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05610_ _01614_ _02096_ _01654_ _02097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_91_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06590_ _02754_ _02834_ _02842_ _00230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_17_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05731__A2 _02167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05541_ _01636_ _02028_ _01417_ _02029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08260_ _03763_ _03828_ _03851_ _03852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09656__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05472_ u_cpu.rf_ram.memory\[4\]\[4\] u_cpu.rf_ram.memory\[5\]\[4\] u_cpu.rf_ram.memory\[6\]\[4\]
+ u_cpu.rf_ram.memory\[7\]\[4\] _01546_ _01550_ _01960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07484__A2 _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07211_ u_cpu.rf_ram.memory\[71\]\[6\] _03186_ _03193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08191_ _03754_ _03755_ _03791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10633__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07142_ _03151_ _00473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08433__A1 _03999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07236__A2 _03206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05247__A1 _01636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08984__A2 _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07073_ _03113_ _00442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_127_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06024_ _02480_ _02481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10783__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08736__A2 _04199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07975_ u_cpu.rf_ram.memory\[116\]\[2\] _03626_ _03629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09714_ _00168_ io_in[4] u_cpu.rf_ram.memory\[47\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05464__B _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10013__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06926_ u_cpu.rf_ram.memory\[58\]\[1\] _03031_ _03033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__04859__I u_cpu.cpu.state.genblk1.misalign_trap_sync_r vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09161__A2 _04449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09645_ _00099_ io_in[4] u_cpu.rf_ram.memory\[42\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06857_ u_cpu.rf_ram.memory\[61\]\[2\] _02992_ _02995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07172__A1 _03169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05808_ _02273_ _02292_ _01402_ _02293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_76_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09576_ _00030_ io_in[4] u_cpu.rf_ram.memory\[82\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06788_ _02754_ _02944_ _02952_ _00318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_42_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05722__A2 _02207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08494__C _03797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10163__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08527_ _04083_ _04084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05739_ _01562_ _02223_ _01565_ _02224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_70_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08458_ u_cpu.cpu.csr_imm _02305_ _03798_ _04014_ _04023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_51_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07409_ _03171_ _03295_ _03302_ _00589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08389_ _03761_ _03860_ _03828_ _03788_ _03800_ _03962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_13_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10420_ _00853_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08424__A1 _01372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07227__A2 _03196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09472__I0 _02573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05238__A1 _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10351_ _00784_ io_in[4] u_cpu.rf_ram.memory\[121\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08975__A2 _04197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10282_ _00715_ io_in[4] u_cpu.rf_ram.memory\[91\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06738__A1 _02738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05410__A1 _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09152__A2 _04439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10506__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07163__A1 _03163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08360__B1 _03779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09679__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08112__B1 _03654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10656__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07466__A2 _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10618_ _01047_ io_in[4] u_cpu.rf_ram.memory\[93\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07218__A2 _03196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05229__A1 _01601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10549_ _00981_ io_in[4] u_cpu.rf_ram.memory\[30\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08718__A2 _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10036__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07256__S _03215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09391__A2 _01377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05401__A1 _01594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07760_ _03355_ _03500_ _03506_ _00737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05284__B _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04972_ _01443_ _01480_ _01481_ _01482_ u_arbiter.o_wb_cpu_adr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_110_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05952__A2 _01403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09143__A2 _04439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10186__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06711_ u_cpu.rf_ram.memory\[68\]\[5\] _02904_ _02910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07691_ _03463_ _00710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07154__A1 _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09430_ _04480_ _04605_ _04611_ _01302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06201__I0 _02587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06642_ _02752_ _02864_ _02871_ _00253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09361_ _02305_ _02344_ _02338_ _04566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_u_scanchain_local.scan_flop\[1\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06573_ _02539_ _02832_ _02833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08312_ _03831_ _03789_ _03892_ _03893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05524_ _01422_ _02002_ _02011_ _02012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_75_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09292_ u_cpu.rf_ram.memory\[86\]\[1\] _04526_ _04528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08654__A1 _02305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07457__A2 _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08243_ _03742_ _03757_ _03836_ _03837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_138_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05455_ _01539_ _01934_ _01943_ _01944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_20_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08406__A1 _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08174_ _03773_ _03755_ _03774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07209__A2 _03186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05386_ u_cpu.rf_ram.memory\[0\]\[3\] u_cpu.rf_ram.memory\[1\]\[3\] u_cpu.rf_ram.memory\[2\]\[3\]
+ u_cpu.rf_ram.memory\[3\]\[3\] _01556_ _01557_ _01875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_118_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07125_ _02959_ _03139_ _03142_ _00465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07056_ _03104_ _00434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06007_ _02459_ _02463_ _02464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05640__A1 _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08489__C _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10529__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[14\]_SI u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07393__A1 _03173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05194__B _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07958_ _03545_ _03616_ _03619_ _00822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09821__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09134__A2 _04429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06909_ _03023_ _00368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07889_ _03581_ _00791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09628_ _00082_ io_in[4] u_cpu.rf_ram.memory\[80\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10679__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07696__A2 _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05251__S0 _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05641__C _01404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09559_ _04484_ _04674_ _04682_ _01360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09971__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07448__A2 _02832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08645__A1 _03547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06120__A2 _02551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10403_ _00836_ io_in[4] u_cpu.rf_ram.memory\[33\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10059__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09070__A1 _04284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10334_ _00767_ io_in[4] u_cpu.rf_ram.memory\[120\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07620__A2 _03422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05631__A1 _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10265_ _00698_ io_in[4] u_cpu.rf_ram.memory\[36\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07076__S _03109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09373__A2 _01393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10196_ _00642_ io_in[4] u_cpu.rf_ram.memory\[127\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09125__A2 _04429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05490__S0 _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07136__A1 _02577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05832__B u_cpu.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05242__S0 _01619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05698__A1 _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05793__S1 _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07439__A2 _03315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08636__A1 _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05123__I _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06111__A2 _02541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05545__S1 _01681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05240_ _01422_ _01721_ _01730_ _01731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__06155__S _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08939__A2 _04322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05870__A1 _02309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05171_ _01609_ _01662_ _01663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07611__A2 _03412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08930_ u_cpu.rf_ram.memory\[28\]\[2\] _04322_ _04325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09844__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08861_ _04280_ _04282_ _04283_ _01061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07375__A1 _03173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07812_ _03353_ _03530_ _03535_ _00760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08792_ u_cpu.rf_ram.memory\[93\]\[4\] _04227_ _04232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10821__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05925__A2 _02356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09116__A2 _04419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07743_ u_cpu.cpu.mem_bytecnt\[1\] _02395_ _00710_ _03497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__05481__S0 _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04955_ u_arbiter.i_wb_cpu_dbus_adr\[10\] _01443_ _01469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07127__A1 _02961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08324__B1 _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08175__I0 u_arbiter.i_wb_cpu_rdt\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09994__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07674_ u_cpu.cpu.state.o_cnt\[2\] u_cpu.cpu.state.o_cnt_r\[3\] _03453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07678__A2 _03454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04886_ u_cpu.cpu.decode.op26 u_cpu.cpu.decode.co_ebreak _01412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05689__A1 _01594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05233__S0 _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06625_ u_cpu.rf_ram.memory\[77\]\[7\] _02854_ _02862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09413_ u_cpu.rf_ram.memory\[27\]\[6\] _04595_ _04602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09344_ u_cpu.rf_ram.memory\[88\]\[0\] _04556_ _04557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06556_ u_cpu.rf_ram.memory\[119\]\[0\] _02823_ _02824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08627__B2 _02445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05507_ _01597_ _01994_ _01995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09275_ _04472_ _04516_ _04518_ _01240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06487_ u_cpu.cpu.state.init_done _01385_ _02433_ _02782_ _02783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__06102__A2 _02541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10201__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05536__S1 _01652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08226_ _02306_ _03798_ _03821_ _03822_ _03823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05438_ _01398_ _01926_ _01927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__04872__I _01397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07850__A2 _03558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05861__A1 _02343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08157_ _03756_ _03757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09052__A1 _04284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05369_ u_cpu.rf_ram.memory\[136\]\[2\] u_cpu.rf_ram.memory\[137\]\[2\] u_cpu.rf_ram.memory\[138\]\[2\]
+ u_cpu.rf_ram.memory\[139\]\[2\] _01680_ _01681_ _01859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_101_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07108_ u_cpu.rf_ram.memory\[141\]\[3\] _03129_ _03133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07602__A2 _03412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08088_ u_arbiter.i_wb_cpu_dbus_dat\[21\] _03683_ _03708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10351__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07039_ _02961_ _03091_ _03095_ _00426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09355__A2 _04556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10050_ _00496_ io_in[4] u_cpu.rf_ram.memory\[71\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05916__A2 _02395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09107__A2 _04419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05472__S0 _01546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07118__A1 _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07669__A2 _03442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10952_ u_cpu.rf_ram_if.wdata1_r\[6\] io_in[4] u_cpu.rf_ram_if.wdata1_r\[5\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07913__I0 _02599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05224__S0 _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10883_ _01312_ io_in[4] u_cpu.rf_ram.memory\[25\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06341__A2 _02686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09717__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09291__A1 _04468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08094__A2 _03653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05527__S1 _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07841__A2 _03541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05852__A1 _01370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09867__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05604__A1 _01589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10317_ _00750_ io_in[4] u_cpu.rf_ram.memory\[34\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_u_scanchain_local.scan_flop\[54\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10844__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09346__A2 _04556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10248_ _00681_ io_in[4] u_cpu.rf_ram.memory\[38\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07357__A1 _03173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10179_ _00625_ io_in[4] u_cpu.rf_ram.memory\[22\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05118__I _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[69\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05463__S0 _01687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07109__A1 _02961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06580__A2 _02834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05215__S0 _01578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06332__A2 _02684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10224__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06410_ _02482_ _02729_ _02730_ _00162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_16_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07390_ u_cpu.rf_ram.memory\[134\]\[6\] _03285_ _03292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__04894__A2 _01388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06341_ _02497_ _02686_ _02690_ _00133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08085__A2 _03683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09060_ _04292_ _04389_ _04395_ _01148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06272_ _02517_ _02641_ _02649_ _00105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07832__A2 _03541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10374__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08011_ u_arbiter.i_wb_cpu_dbus_dat\[1\] _02774_ _02781_ _03651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05843__A1 _02309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05223_ _01589_ _01713_ _01714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09034__A1 _04284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05154_ _01544_ _01646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07596__A1 _03357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06399__A2 _02718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05085_ _01543_ _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09962_ _00416_ io_in[4] u_cpu.rf_ram.memory\[53\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08913_ u_cpu.rf_ram.memory\[96\]\[5\] _04309_ _04315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09337__A2 _04546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09893_ _00347_ io_in[4] u_cpu.rf_ram.memory\[61\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08844_ _03543_ _04271_ _04273_ _01054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08775_ _04222_ _01036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05987_ u_arbiter.i_wb_cpu_ibus_adr\[0\] u_cpu.cpu.ctrl.pc_plus_4_cy_r _02450_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06571__A2 _02823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07726_ u_cpu.rf_ram.memory\[90\]\[7\] _03475_ _03483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04938_ _01431_ _01455_ _01456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08848__A1 _03547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05206__S0 _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07657_ u_cpu.rf_ram.memory\[36\]\[1\] _03442_ _03444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04869_ _01393_ _01394_ _01387_ _01368_ _01395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__06323__A2 _02673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07520__A1 _03353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06608_ _02754_ _02844_ _02852_ _00238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07588_ _03349_ _03402_ _03405_ _00665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_90_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10717__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06539_ u_cpu.rf_ram.memory\[40\]\[1\] _02812_ _02814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09327_ _04468_ _04546_ _04547_ _01263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09273__A1 _04468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06087__A1 _02492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09258_ u_cpu.rf_ram.memory\[85\]\[2\] _04506_ _04509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07823__A2 _03541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05834__A1 _02311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08209_ _03765_ _03778_ _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_09189_ u_cpu.rf_ram.memory\[69\]\[7\] _04459_ _04467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10867__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05647__B _01417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10102_ _00548_ io_in[4] u_cpu.rf_ram.memory\[137\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09328__A2 _04546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11082_ _11082_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__05693__S0 _01646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05366__C _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07339__A1 _03173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10033_ _00479_ io_in[4] u_cpu.rf_ram.memory\[72\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08000__A2 _03636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06011__A1 _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06562__A2 _02823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10247__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08839__A1 _02539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07153__I _02481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09500__A2 _04644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10935_ u_cpu.rf_ram_if.wdata0_r\[2\] io_in[4] u_cpu.rf_ram_if.wdata0_r\[1\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06314__A2 _02673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05373__I0 u_cpu.rf_ram.memory\[128\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10866_ _01295_ io_in[4] u_cpu.rf_ram.memory\[27\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10397__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08067__A2 _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10797_ _01226_ io_in[4] u_cpu.rf_ram.memory\[10\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06078__A1 u_cpu.cpu.immdec.imm11_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07814__A2 _03530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09016__A1 _04284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07578__A1 _03357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09319__A2 _04536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05684__S0 _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05910_ _01372_ _02313_ _02391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06890_ _02953_ _03012_ _03013_ _00359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_79_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07264__S _03215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05841_ _02319_ _02324_ _02306_ _02325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07750__A1 _03343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05772_ u_cpu.rf_ram.memory\[104\]\[7\] u_cpu.rf_ram.memory\[105\]\[7\] u_cpu.rf_ram.memory\[106\]\[7\]
+ u_cpu.rf_ram.memory\[107\]\[7\] _01615_ _01616_ _02257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_48_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08560_ u_cpu.rf_ram.memory\[31\]\[7\] _04094_ _04102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07511_ u_cpu.rf_ram.memory\[128\]\[0\] _03362_ _03363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08491_ _03849_ _03897_ _04053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06305__A2 _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07502__A1 _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07442_ u_cpu.rf_ram.memory\[131\]\[5\] _03315_ _03321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04867__A2 u_cpu.cpu.state.genblk1.misalign_trap_sync_r vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07373_ _03171_ _03275_ _03282_ _00573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09255__A1 _04468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08058__A2 _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06069__A1 _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09112_ _04290_ _04419_ _04424_ _01171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06324_ _02507_ _02673_ _02679_ _00127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07805__A2 _03530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09043_ u_cpu.rf_ram.memory\[104\]\[6\] _04379_ _04386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05816__A1 _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06255_ _02638_ _02639_ _02640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05206_ u_cpu.rf_ram.memory\[12\]\[1\] u_cpu.rf_ram.memory\[13\]\[1\] u_cpu.rf_ram.memory\[14\]\[1\]
+ u_cpu.rf_ram.memory\[15\]\[1\] _01556_ _01557_ _01697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09558__A2 _04674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06186_ _02596_ u_cpu.rf_ram.memory\[1\]\[6\] _02578_ _02597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05137_ _01613_ _01618_ _01622_ _01627_ _01628_ _01629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_143_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08230__A2 _03755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06241__A1 _02492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05675__S0 _01619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05068_ u_cpu.rf_ram.memory\[4\]\[0\] u_cpu.rf_ram.memory\[5\]\[0\] u_cpu.rf_ram.memory\[6\]\[0\]
+ u_cpu.rf_ram.memory\[7\]\[0\] _01546_ _01550_ _01560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09945_ _00399_ io_in[4] u_cpu.rf_ram.memory\[55\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06792__A2 _02955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09876_ _00330_ io_in[4] u_cpu.rf_ram.memory\[63\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05427__S0 _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08827_ _03778_ _03780_ _04259_ _03742_ _04260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_38_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06544__A2 _02812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07741__A1 _02313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08758_ _04213_ _01028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_73_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07709_ _03359_ _03465_ _03473_ _00718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08297__A2 _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08689_ u_cpu.cpu.ctrl.o_ibus_adr\[15\] _04173_ _04157_ u_cpu.cpu.ctrl.o_ibus_adr\[16\]
+ _04174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10720_ _01149_ io_in[4] u_cpu.rf_ram.memory\[99\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10651_ _01080_ io_in[4] u_cpu.rf_ram.memory\[96\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08018__B _02774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10582_ _01012_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05807__A1 _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09549__A2 _04674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08221__A2 _03802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05666__S0 _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05096__C _01426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07980__A1 _03549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06783__A2 _02944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09905__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11065_ _11065_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_122_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05418__S0 _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10016_ _00462_ io_in[4] u_cpu.rf_ram.memory\[141\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08524__A3 u_cpu.cpu.genblk3.csr.i_mtip vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05824__C _01374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06535__A2 _02810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08780__I0 _02599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08288__A2 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06299__A1 _02492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10918_ _01347_ io_in[4] u_cpu.rf_ram.memory\[89\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10849_ _01278_ io_in[4] u_cpu.rf_ram.memory\[88\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_u_scanchain_local.scan_flop\[40\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05131__I _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08460__A2 _03988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06040_ _02478_ u_cpu.rf_ram_if.wdata1_r\[3\] _02494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_132_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xu_scanchain_local.output_buffers\[2\] u_scanchain_local.data_out_i u_scanchain_local.data_out
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_114_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08212__A2 _03809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10412__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06223__A1 _02502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09474__S _04634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05657__S0 _01546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07991_ u_cpu.rf_ram.memory\[33\]\[1\] _03636_ _03638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09585__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06774__A2 _02944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09730_ _00184_ io_in[4] u_cpu.rf_ram.memory\[4\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06942_ u_cpu.rf_ram.memory\[57\]\[0\] _03041_ _03042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05409__S0 _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09661_ _00115_ io_in[4] u_cpu.rf_ram.memory\[45\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10562__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06873_ u_cpu.rf_ram.memory\[60\]\[1\] _03002_ _03004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07723__A1 _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05329__A3 _01799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06526__A2 _02801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08612_ _04128_ _00967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05824_ _02306_ u_cpu.cpu.bufreg.i_sh_signed _02307_ _01374_ _02308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_82_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09592_ _00046_ io_in[4] u_cpu.rf_ram.memory\[81\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08543_ _03555_ _04084_ _04092_ _00934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05755_ _01636_ _02239_ _02240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05686_ u_cpu.rf_ram.memory\[100\]\[6\] u_cpu.rf_ram.memory\[101\]\[6\] u_cpu.rf_ram.memory\[102\]\[6\]
+ u_cpu.rf_ram.memory\[103\]\[6\] _01577_ _01549_ _02172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08474_ u_arbiter.i_wb_cpu_rdt\[16\] u_arbiter.i_wb_cpu_rdt\[0\] _01436_ _04037_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_126_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07425_ _03169_ _03305_ _03311_ _00596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09228__A1 _04478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07356_ u_cpu.rf_ram.memory\[136\]\[7\] _03265_ _03273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06307_ _02512_ _02662_ _02669_ _00120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07287_ _03234_ _03235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07677__B _01429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09026_ _04294_ _04369_ _04376_ _01133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06238_ u_cpu.rf_ram.memory\[78\]\[1\] _02628_ _02630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09928__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10092__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06169_ _02583_ _02584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_46_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07262__I0 _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05648__S0 _01578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10905__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07962__A1 _03549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06765__A2 _02934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09928_ _00382_ io_in[4] u_cpu.rf_ram.memory\[58\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09859_ _00313_ io_in[4] u_cpu.rf_ram.memory\[64\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07190__A2 _03176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05660__B _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[63\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10703_ _01132_ io_in[4] u_cpu.rf_ram.memory\[103\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10634_ _01063_ io_in[4] u_cpu.rf_ram.memory\[94\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10565_ _00995_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10435__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05256__A2 _01746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10496_ _00929_ io_in[4] u_cpu.rf_ram.memory\[32\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[33\] u_arbiter.i_wb_cpu_rdt\[30\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[27\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_64_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05008__A2 _01442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05639__S0 _01687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10585__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06756__A2 _02934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11048_ _11048_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07705__A1 _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06508__A2 _02791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08753__I0 _02584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07181__A2 _03176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05811__S0 _01680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09458__A1 _04472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05540_ u_cpu.rf_ram.memory\[76\]\[4\] u_cpu.rf_ram.memory\[77\]\[4\] u_cpu.rf_ram.memory\[78\]\[4\]
+ u_cpu.rf_ram.memory\[79\]\[4\] _01577_ _01549_ _02028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_17_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05471_ _01554_ _01958_ _01417_ _01959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_32_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07210_ _03169_ _03186_ _03192_ _00500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08190_ _03785_ _03787_ _03789_ _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_07141_ _02584_ u_cpu.rf_ram.memory\[13\]\[2\] _03148_ _03151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_9_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05247__A2 _01737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06444__A1 _02750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07072_ _02587_ u_cpu.rf_ram.memory\[15\]\[3\] _03109_ _03113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05729__C _01404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10928__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06023_ u_cpu.rf_ram_if.wdata0_r\[0\] _02460_ _02479_ _02480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_114_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08197__A1 u_arbiter.i_wb_cpu_ack vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07944__A1 _03549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06747__A2 _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07974_ _03543_ _03626_ _03628_ _00829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09713_ _00167_ io_in[4] u_cpu.rf_ram.memory\[47\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06925_ _02953_ _03031_ _03032_ _00375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09644_ _00098_ io_in[4] u_cpu.rf_ram.memory\[42\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06856_ _02957_ _02992_ _02994_ _00344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07172__A2 _03159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10308__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05807_ _01539_ _02282_ _02291_ _02292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__05802__S0 _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09575_ _00029_ io_in[4] u_cpu.rf_ram.memory\[82\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06787_ u_cpu.rf_ram.memory\[64\]\[7\] _02944_ _02952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08526_ _02612_ _02639_ _04083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05480__B _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04930__A1 u_arbiter.i_wb_cpu_dbus_adr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05738_ u_cpu.rf_ram.memory\[0\]\[7\] u_cpu.rf_ram.memory\[1\]\[7\] u_cpu.rf_ram.memory\[2\]\[7\]
+ u_cpu.rf_ram.memory\[3\]\[7\] _01556_ _01557_ _02223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_70_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09600__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08457_ u_cpu.cpu.immdec.imm19_12_20\[3\] _04016_ _04022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08672__A2 _04155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05669_ _01601_ _02154_ _01605_ _02155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10458__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07408_ u_cpu.rf_ram.memory\[133\]\[6\] _03295_ _03302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08388_ _03756_ _03810_ _03958_ _03960_ _03961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_11_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07339_ _03173_ _03255_ _03263_ _00558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09750__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08424__A2 _02313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05238__A2 _01728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06435__A1 _02744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10350_ _00783_ io_in[4] u_cpu.rf_ram.memory\[121\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06986__A2 _03061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09009_ u_cpu.rf_ram.memory\[102\]\[7\] _04359_ _04367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10281_ _00714_ io_in[4] u_cpu.rf_ram.memory\[91\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06738__A2 _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05410__A2 _01898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08360__A1 _03741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07163__A2 _03159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08360__B2 _03935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06486__B _02781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08112__A1 u_arbiter.i_wb_cpu_rdt\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07161__I _02491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05316__I3 u_cpu.rf_ram.memory\[59\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06674__A1 _02748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10617_ _01046_ io_in[4] u_cpu.rf_ram.memory\[93\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06426__A1 _02469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05229__A2 _01719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10548_ _00980_ io_in[4] u_cpu.rf_ram.memory\[30\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__04988__A1 _01445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10479_ _00912_ io_in[4] u_cpu.cpu.immdec.imm30_25\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08179__A1 _03776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07926__A1 _03549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06729__A2 _02914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05401__A2 _01889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04971_ u_arbiter.i_wb_cpu_dbus_adr\[13\] _01442_ _01482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06710_ _02748_ _02904_ _02909_ _00283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_49_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07690_ _01429_ u_cpu.cpu.state.o_cnt_r\[2\] _03463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_92_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09623__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08351__A1 _03776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07154__A2 _02810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05165__A1 _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06641_ u_cpu.rf_ram.memory\[74\]\[6\] _02864_ _02871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06901__A2 _03012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09360_ _02311_ _01386_ _04565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10600__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06572_ _02457_ _02471_ _02832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08103__A1 _02781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08311_ _03785_ _03787_ _03892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_75_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05523_ _02004_ _02006_ _02008_ _02010_ _01607_ _02011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_09291_ _04468_ _04526_ _04527_ _01247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09773__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08654__A2 _02448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08242_ _03741_ _03818_ _03836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05454_ _01936_ _01938_ _01940_ _01942_ _01568_ _01943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_119_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10750__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05385_ _01554_ _01873_ _01874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08173_ _03772_ _03773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07124_ u_cpu.rf_ram.memory\[140\]\[2\] _03139_ _03142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08831__S _03797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06968__A2 _03051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07055_ _02587_ u_cpu.rf_ram.memory\[9\]\[3\] _03100_ _03104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_134_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06006_ _01386_ _02462_ _02463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05640__A2 _02126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08965__I0 u_arbiter.i_wb_cpu_rdt\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05475__B _01565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07393__A2 _03285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10130__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07957_ u_cpu.rf_ram.memory\[115\]\[2\] _03616_ _03619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06908_ _02581_ u_cpu.rf_ram.memory\[5\]\[1\] _03021_ _03023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07888_ _02587_ u_cpu.rf_ram.memory\[8\]\[3\] _03577_ _03581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08342__A1 _03866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09627_ _00081_ io_in[4] u_cpu.rf_ram.memory\[7\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06839_ u_cpu.rf_ram.memory\[62\]\[2\] _02982_ _02985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08893__A2 _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10280__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05251__S1 _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09558_ u_cpu.rf_ram.memory\[23\]\[7\] _04674_ _04682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08509_ _01437_ _03668_ _04069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09489_ _04643_ _04644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08645__A2 _04145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06656__A1 _02748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10402_ _00835_ io_in[4] u_cpu.rf_ram.memory\[116\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09070__A2 _04399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10333_ _00766_ io_in[4] u_cpu.rf_ram.memory\[120\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05631__A2 _02108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10264_ _00697_ io_in[4] u_cpu.rf_ram.memory\[36\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10195_ _00641_ io_in[4] u_cpu.rf_ram.memory\[127\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09646__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07384__A2 _03285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05490__S1 _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08188__S _01435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10623__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07136__A2 _02660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06195__I0 _02573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09796__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05242__S1 _01620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10773__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08097__B1 _03654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08636__A2 _02625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10003__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05170_ u_cpu.rf_ram.memory\[80\]\[0\] u_cpu.rf_ram.memory\[81\]\[0\] u_cpu.rf_ram.memory\[82\]\[0\]
+ u_cpu.rf_ram.memory\[83\]\[0\] _01545_ _01642_ _01662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_7_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05870__A2 _02325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09061__A2 _04389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10153__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08947__I0 u_arbiter.i_wb_cpu_rdt\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05295__B _01417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08860_ u_cpu.rf_ram.memory\[94\]\[0\] _04282_ _04283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09482__S _04634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07375__A2 _03275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07811_ u_cpu.rf_ram.memory\[117\]\[4\] _03530_ _03535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08791_ _03547_ _04227_ _04231_ _01043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07742_ _03486_ _03496_ _00729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04954_ _01445_ _01467_ _01468_ u_arbiter.o_wb_cpu_adr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05481__S1 _01574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08324__A1 _03744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07127__A2 _03139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08324__B2 _03890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05138__A1 _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07673_ _03452_ _00703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06186__I0 _02596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08875__A2 _04282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04885_ _01410_ _01376_ _01411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09412_ _04480_ _04595_ _04601_ _01294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05233__S1 _01616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06624_ _02752_ _02854_ _02861_ _00245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_92_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06886__A1 _02969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09343_ _04555_ _04556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06555_ _02822_ _02823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05506_ u_cpu.rf_ram.memory\[108\]\[4\] u_cpu.rf_ram.memory\[109\]\[4\] u_cpu.rf_ram.memory\[110\]\[4\]
+ u_cpu.rf_ram.memory\[111\]\[4\] _01598_ _01573_ _01994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06638__A1 _02748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09274_ u_cpu.rf_ram.memory\[110\]\[1\] _04516_ _04518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06486_ _01373_ _02780_ _02781_ _01375_ _02782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_21_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08225_ _03754_ _03778_ _03782_ _03759_ _03797_ _03822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_05437_ u_cpu.rf_ram.memory\[92\]\[3\] u_cpu.rf_ram.memory\[93\]\[3\] u_cpu.rf_ram.memory\[94\]\[3\]
+ u_cpu.rf_ram.memory\[95\]\[3\] _01610_ _01611_ _01926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_21_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08156_ u_arbiter.i_wb_cpu_rdt\[6\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[6\]
+ _01435_ _03756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__05861__A2 u_cpu.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05368_ _01838_ _01857_ _01402_ _01858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09052__A2 _04389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07107_ _02959_ _03129_ _03132_ _00457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07685__B _02433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08087_ _03706_ _03707_ _00863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05299_ _01562_ _01788_ _01565_ _01789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09669__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06810__A1 u_cpu.rf_ram.memory\[29\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07038_ u_cpu.rf_ram.memory\[52\]\[3\] _03091_ _03095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10646__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08563__A1 _02433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07366__A2 _03275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07905__S _03586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08989_ u_cpu.rf_ram.memory\[101\]\[6\] _04349_ _04356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05472__S1 _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08315__A1 _03776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07118__A2 _02832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09191__I _02481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10796__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10951_ u_cpu.rf_ram_if.wdata1_r\[5\] io_in[4] u_cpu.rf_ram_if.wdata1_r\[4\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05652__C _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08866__A2 _04282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05224__S1 _01548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10882_ _01311_ io_in[4] u_cpu.rf_ram.memory\[25\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10026__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09291__A2 _04526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06055__I _02506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10176__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09043__A2 _04379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08251__B1 _03801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10316_ _00749_ io_in[4] u_cpu.rf_ram.memory\[34\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05604__A2 _02090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06801__A1 u_cpu.rf_ram.memory\[29\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10247_ _00680_ io_in[4] u_cpu.rf_ram.memory\[38\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07357__A2 _03265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05368__A1 _01838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10178_ _00624_ io_in[4] u_cpu.rf_ram.memory\[22\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05463__S1 _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08306__A1 _03555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07109__A2 _03129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06868__A1 _02969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05215__S1 _01580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05134__I _01564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06340_ u_cpu.rf_ram.memory\[51\]\[3\] _02686_ _02690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06166__S _02578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09282__A2 _04516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10519__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06271_ u_cpu.rf_ram.memory\[42\]\[7\] _02641_ _02649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06096__A2 _02530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07293__A1 _03163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08010_ _03648_ _03649_ _03650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05222_ u_cpu.rf_ram.memory\[52\]\[1\] u_cpu.rf_ram.memory\[53\]\[1\] u_cpu.rf_ram.memory\[54\]\[1\]
+ u_cpu.rf_ram.memory\[55\]\[1\] _01590_ _01591_ _01713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09811__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09034__A2 _04379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05153_ _01540_ _01645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07045__A1 _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10669__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07596__A2 _03402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08793__A1 _03549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09961_ _00415_ io_in[4] u_cpu.rf_ram.memory\[53\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05084_ _01570_ _01575_ _01576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05151__S0 _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08912_ _04290_ _04309_ _04314_ _01081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09961__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09892_ _00346_ io_in[4] u_cpu.rf_ram.memory\[61\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07348__A2 _03265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08843_ u_cpu.rf_ram.memory\[97\]\[1\] _04271_ _04273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05359__A1 _01667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05753__B _01564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08774_ _02590_ u_cpu.rf_ram.memory\[2\]\[4\] _04217_ _04222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_100_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05986_ _02446_ _02404_ _02449_ _00024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07725_ _03357_ _03475_ _03482_ _00725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04937_ u_cpu.cpu.ctrl.o_ibus_adr\[6\] u_cpu.cpu.ctrl.o_ibus_adr\[5\] _01451_ _01455_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_66_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08848__A2 _04271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10049__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05206__S1 _01557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07656_ _03343_ _03442_ _03443_ _00695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_04868_ u_cpu.cpu.decode.op21 _01380_ _01394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_26_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07520__A2 _03362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06607_ u_cpu.rf_ram.memory\[139\]\[7\] _02844_ _02852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07587_ u_cpu.rf_ram.memory\[124\]\[2\] _03402_ _03405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09326_ u_cpu.rf_ram.memory\[87\]\[0\] _04546_ _04547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06538_ _02738_ _02812_ _02813_ _00207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10199__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09273__A2 _04516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06087__A2 _02530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09257_ _04472_ _04506_ _04508_ _01232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06469_ u_arbiter.i_wb_cpu_ack _01431_ _02766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08208_ _03798_ _03805_ _03806_ _00885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05834__A2 u_cpu.cpu.immdec.imm31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09188_ _04294_ _04459_ _04466_ _01205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09025__A2 _04369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08139_ _03555_ _03731_ _03739_ _00883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07587__A2 _03402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05142__S0 _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10101_ _00547_ io_in[4] u_cpu.rf_ram.memory\[137\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11081_ _11081_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__05693__S1 _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[1\]_D u_cpu.cpu.genblk3.csr.i_mtip vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07339__A2 _03255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10032_ _00478_ io_in[4] u_cpu.rf_ram.memory\[13\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08839__A2 _04197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10934_ u_cpu.rf_ram_if.wdata0_r\[1\] io_in[4] u_cpu.rf_ram_if.wdata0_r\[0\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07511__A2 _03362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05522__A1 _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10865_ _01294_ io_in[4] u_cpu.rf_ram.memory\[27\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09834__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09264__A2 _04506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10796_ _01225_ io_in[4] u_cpu.rf_ram.memory\[10\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[63\] u_scanchain_local.module_data_in\[62\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[25\] u_scanchain_local.clk u_scanchain_local.module_data_in\[63\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__07275__A1 _03163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10811__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09016__A2 _04369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07027__A1 _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09984__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07578__A2 _03392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05133__S0 _01623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06250__A2 _02628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05684__S1 _01616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05840_ _02320_ _02322_ _02323_ _02324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_82_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07750__A2 _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05771_ _01597_ _02255_ _02256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07510_ _03361_ _03362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08490_ _03782_ _04051_ _04052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_63_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07502__A2 _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10341__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07441_ _03167_ _03315_ _03320_ _00603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05513__A1 _01601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07372_ u_cpu.rf_ram.memory\[135\]\[6\] _03275_ _03282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09255__A2 _04506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09111_ u_cpu.rf_ram.memory\[106\]\[4\] _04419_ _04424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06323_ u_cpu.rf_ram.memory\[44\]\[5\] _02673_ _02679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06069__A2 _02517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10491__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09042_ _04292_ _04379_ _04385_ _01140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05816__A2 _02300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06254_ u_cpu.cpu.immdec.imm11_7\[2\] _02526_ _02574_ _02639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__09007__A2 _04359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05205_ _01542_ _01695_ _01696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05748__B _01417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06185_ _02595_ _02596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07569__A2 _03392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05136_ _01567_ _01628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05067_ _01554_ _01558_ _01417_ _01559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09944_ _00398_ io_in[4] u_cpu.rf_ram.memory\[56\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06241__A2 _02628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05675__S1 _01620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08518__A1 _03835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09875_ _00329_ io_in[4] u_cpu.rf_ram.memory\[63\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09707__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05427__S1 _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08826_ _03755_ _03786_ _04256_ _03851_ _04259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08757_ _02590_ u_cpu.rf_ram.memory\[3\]\[4\] _04208_ _04213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_45_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05969_ _02432_ _02435_ _01445_ u_arbiter.o_wb_cpu_cyc vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07708_ u_cpu.rf_ram.memory\[91\]\[7\] _03465_ _03473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08688_ _04154_ _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09857__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09494__A2 _04644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07639_ u_cpu.rf_ram.memory\[37\]\[1\] _03432_ _03434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05504__A1 _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[53\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10650_ _01079_ io_in[4] u_cpu.rf_ram.memory\[96\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10834__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09309_ _04468_ _04536_ _04537_ _01255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10581_ _01011_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05807__A2 _02282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[68\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07009__A1 _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08034__B _03648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05377__C _01404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10214__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05666__S1 _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08509__A1 _01437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07980__A2 _03626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11064_ _11064_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_122_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09182__A1 _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10015_ _00461_ io_in[4] u_cpu.rf_ram.memory\[141\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05418__S1 _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07164__I _02496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10364__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10917_ _01346_ io_in[4] u_cpu.rf_ram.memory\[89\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06299__A2 _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07496__A1 _03351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10848_ _01277_ io_in[4] u_cpu.rf_ram.memory\[88\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_u_scanchain_local.scan_flop\[34\]_D u_arbiter.i_wb_cpu_rdt\[31\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07248__A1 _03171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10779_ _01208_ io_in[4] u_cpu.rf_ram.memory\[84\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07799__A2 _03520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08996__A1 _04280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05568__B _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08748__A1 _02577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06223__A2 _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05657__S1 _01574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07990_ _03539_ _03636_ _03637_ _00836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07971__A2 _03626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06941_ _03040_ _03041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10707__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05982__A1 u_arbiter.i_wb_cpu_ibus_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09173__A1 _02524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05409__S1 _01616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09660_ _00114_ io_in[4] u_cpu.rf_ram.memory\[45\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06872_ _02953_ _03002_ _03003_ _00351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07723__A2 _03475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08920__A1 _03991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08611_ u_arbiter.i_wb_cpu_dbus_adr\[26\] u_arbiter.i_wb_cpu_dbus_adr\[25\] _04115_
+ _04128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05823_ _01409_ _02307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09591_ _00045_ io_in[4] u_cpu.rf_ram.memory\[81\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08542_ u_cpu.rf_ram.memory\[32\]\[7\] _04084_ _04092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10857__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05754_ u_cpu.rf_ram.memory\[60\]\[7\] u_cpu.rf_ram.memory\[61\]\[7\] u_cpu.rf_ram.memory\[62\]\[7\]
+ u_cpu.rf_ram.memory\[63\]\[7\] _01598_ _01573_ _02239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_82_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07487__A1 _03343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08473_ _01390_ _04016_ _04035_ _04036_ _00920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_39_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05685_ _01594_ _02170_ _01416_ _02171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08684__B1 _04157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07424_ u_cpu.rf_ram.memory\[132\]\[5\] _03305_ _03311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_u_scanchain_local.scan_flop\[25\]_D u_arbiter.i_wb_cpu_rdt\[22\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09228__A2 _04487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07355_ _03171_ _03265_ _03272_ _00565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06306_ u_cpu.rf_ram.memory\[45\]\[6\] _02662_ _02669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05345__S0 _01623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07286_ _02602_ _02639_ _03234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09025_ u_cpu.rf_ram.memory\[103\]\[6\] _04369_ _04376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06237_ _02482_ _02628_ _02629_ _00090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10237__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08739__A1 _03547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06168_ u_cpu.rf_ram_if.wdata0_r\[2\] u_cpu.rf_ram_if.wdata1_r\[2\] _02478_ _02583_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06214__A2 _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05119_ _01548_ _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07411__A1 _03173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05648__S1 _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06099_ _02475_ _02539_ _02540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07962__A2 _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10387__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09927_ _00381_ io_in[4] u_cpu.rf_ram.memory\[58\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05973__A1 _01374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09164__A1 _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09858_ _00312_ io_in[4] u_cpu.rf_ram.memory\[64\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07714__A2 _03475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07913__S _03586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08809_ _03780_ _04243_ _04244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09789_ _00243_ io_in[4] u_cpu.rf_ram.memory\[77\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09467__A2 _04625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10702_ _01131_ io_in[4] u_cpu.rf_ram.memory\[103\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06150__A1 _02507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[16\]_D u_arbiter.i_wb_cpu_rdt\[13\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09219__A2 _04487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10633_ _01062_ io_in[4] u_cpu.rf_ram.memory\[94\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08978__A1 _04280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10564_ _00994_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05336__S0 _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07650__A1 _03357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10495_ _00928_ io_in[4] u_cpu.rf_ram.memory\[32\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[26\] u_arbiter.i_wb_cpu_rdt\[23\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[20\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__05639__S1 _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07953__A2 _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09155__A1 _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11047_ _11047_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_77_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07705__A2 _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08363__C1 _03935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05811__S1 _01681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09458__A2 _04625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08666__B1 _04157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08130__A2 _03731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05470_ u_cpu.rf_ram.memory\[12\]\[4\] u_cpu.rf_ram.memory\[13\]\[4\] u_cpu.rf_ram.memory\[14\]\[4\]
+ u_cpu.rf_ram.memory\[15\]\[4\] _01556_ _01557_ _01958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_20_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07140_ _03150_ _00472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06174__S _02578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07071_ _03112_ _00441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06444__A2 _02740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06022_ u_cpu.rf_ram_if.wdata1_r\[0\] _02478_ _02479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_127_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08197__A2 _01431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07944__A2 _03606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07973_ u_cpu.rf_ram.memory\[116\]\[1\] _03626_ _03628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05955__A1 _01403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09146__A1 _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09712_ _00166_ io_in[4] u_cpu.rf_ram.memory\[47\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_101_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06924_ u_cpu.rf_ram.memory\[58\]\[0\] _03031_ _03032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09643_ _00097_ io_in[4] u_cpu.rf_ram.memory\[78\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06855_ u_cpu.rf_ram.memory\[61\]\[1\] _02992_ _02994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05806_ _02284_ _02286_ _02288_ _02290_ _01568_ _02291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_27_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09574_ _00028_ io_in[4] u_cpu.rf_ram.memory\[82\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05802__S1 _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06786_ _02752_ _02944_ _02951_ _00317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09449__A2 _04615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08525_ _04080_ _04081_ _04082_ _00926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05737_ _01554_ _02221_ _02222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04930__A2 _01443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08121__A2 _03678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08456_ _04020_ _04016_ _04021_ _03840_ _00918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_23_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08564__S _02445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05668_ u_cpu.rf_ram.memory\[56\]\[6\] u_cpu.rf_ram.memory\[57\]\[6\] u_cpu.rf_ram.memory\[58\]\[6\]
+ u_cpu.rf_ram.memory\[59\]\[6\] _01602_ _01579_ _02154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06132__A1 _02512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05052__I _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07407_ _03169_ _03295_ _03301_ _00588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07880__A1 _03555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08387_ _03773_ _03959_ _03960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05599_ _01636_ _02085_ _02086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04891__I _01416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07338_ u_cpu.rf_ram.memory\[49\]\[7\] _03255_ _03263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07632__A1 _03357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06435__A2 _02740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07269_ _03224_ _03225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09008_ _04294_ _04359_ _04366_ _01125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10280_ _00713_ io_in[4] u_cpu.rf_ram.memory\[91\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07935__A2 _03606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05946__A1 _02320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09137__A1 _02475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[30\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07699__A1 _03349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08360__A2 _03778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06486__C _01375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08112__A2 _03653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10402__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08474__S _01436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09575__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06674__A2 _02884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10616_ _01045_ io_in[4] u_cpu.rf_ram.memory\[93\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10552__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10455__D _00888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06426__A2 _02684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10547_ _00979_ io_in[4] u_cpu.rf_ram.memory\[30\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10478_ _00911_ io_in[4] u_cpu.cpu.immdec.imm30_25\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08179__A2 _03778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07926__A2 _03596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05937__A1 _02320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09128__A1 _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04970_ u_cpu.cpu.ctrl.o_ibus_adr\[13\] u_cpu.cpu.ctrl.o_ibus_adr\[12\] _01476_ _01481_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_49_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08351__A2 _03923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06640_ _02750_ _02864_ _02870_ _00252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05581__B _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05165__A2 _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06362__A1 _02502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06571_ _02754_ _02823_ _02831_ _00222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09918__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08310_ _03745_ _03788_ _03891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08103__A2 _03648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10082__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05522_ _01614_ _02009_ _01654_ _02010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09290_ u_cpu.rf_ram.memory\[86\]\[0\] _04526_ _04527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06114__A1 _02512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08241_ _03751_ _03803_ _03835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07862__A1 _03555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05453_ _01636_ _01941_ _01417_ _01942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06665__A2 _02884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08172_ u_arbiter.i_wb_cpu_rdt\[0\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[0\]
+ _01435_ _03772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05384_ u_cpu.rf_ram.memory\[4\]\[3\] u_cpu.rf_ram.memory\[5\]\[3\] u_cpu.rf_ram.memory\[6\]\[3\]
+ u_cpu.rf_ram.memory\[7\]\[3\] _01546_ _01550_ _01873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07123_ _02957_ _03139_ _03141_ _00464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06417__A2 _02729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07614__A1 _03357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07054_ _03103_ _00433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07090__A2 _03119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06005_ _02460_ _01412_ _02461_ _02462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09367__A1 _04568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07917__A2 _03596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[53\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05928__A1 _01374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09119__A1 _02706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07956_ _03543_ _03616_ _03618_ _00821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06907_ _03022_ _00367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07887_ _03580_ _00790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_46_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10425__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09626_ _00080_ io_in[4] u_cpu.rf_ram.memory\[7\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06838_ _02957_ _02982_ _02984_ _00336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09598__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09557_ _04482_ _04674_ _04681_ _01359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06769_ u_cpu.rf_ram.memory\[65\]\[7\] _02934_ _02942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08508_ _03849_ _04067_ _04068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09488_ _02469_ _04197_ _04643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10575__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08439_ _03763_ _03778_ _03779_ _03744_ _03851_ _04008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__06656__A2 _02874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10401_ _00834_ io_in[4] u_cpu.rf_ram.memory\[116\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10332_ _00765_ io_in[4] u_cpu.rf_ram.memory\[120\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10263_ _00696_ io_in[4] u_cpu.rf_ram.memory\[36\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05631__A3 _02117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10194_ _00640_ io_in[4] u_cpu.rf_ram.memory\[127\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05919__A1 u_cpu.cpu.decode.opcode\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08333__A2 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06895__A2 _03012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10918__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08097__A1 u_arbiter.i_wb_cpu_rdt\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07844__A1 _03555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06647__A2 _02874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06452__S _02756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09349__A1 _04474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07810_ _03351_ _03530_ _03534_ _00759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10448__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08790_ u_cpu.rf_ram.memory\[93\]\[3\] _04227_ _04231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07741_ _02313_ _03495_ _00703_ _01374_ _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_04953_ u_arbiter.i_wb_cpu_dbus_adr\[9\] _01457_ _01468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09740__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09521__A1 _04482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08324__A2 _03786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07672_ _01428_ _03451_ _03452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_04884_ _01408_ _01409_ _01410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06335__A1 _02482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09411_ u_cpu.rf_ram.memory\[27\]\[5\] _04595_ _04601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06623_ u_cpu.rf_ram.memory\[77\]\[6\] _02854_ _02861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10598__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06886__A2 _03002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09342_ _02475_ _02810_ _04555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06554_ _02602_ _02821_ _02822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09890__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05505_ _01539_ _01964_ _01973_ _01992_ _01993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__07835__A1 _03549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09273_ _04468_ _04516_ _04517_ _01239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06638__A2 _02864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06485_ u_arbiter.i_wb_cpu_ack _01442_ _02781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08224_ _03791_ _03820_ _03821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05436_ _01422_ _01915_ _01924_ _01925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_20_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08155_ u_arbiter.i_wb_cpu_rdt\[1\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\]
+ _01435_ _03755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05861__A3 _01411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05367_ _01539_ _01847_ _01856_ _01857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_07106_ u_cpu.rf_ram.memory\[141\]\[2\] _03129_ _03132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08260__A1 _03763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08086_ u_arbiter.i_wb_cpu_rdt\[19\] _03669_ _03678_ u_arbiter.i_wb_cpu_dbus_dat\[19\]
+ _03707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05298_ u_cpu.rf_ram.memory\[0\]\[2\] u_cpu.rf_ram.memory\[1\]\[2\] u_cpu.rf_ram.memory\[2\]\[2\]
+ u_cpu.rf_ram.memory\[3\]\[2\] _01556_ _01557_ _01788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07685__C _01429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05074__A1 _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07037_ _02959_ _03091_ _03094_ _00425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06810__A2 _02955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08012__A1 u_arbiter.i_wb_cpu_ack vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08988_ _04292_ _04349_ _04355_ _01116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07939_ u_cpu.rf_ram.memory\[122\]\[2\] _03606_ _03609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08315__A2 _03768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10950_ u_cpu.rf_ram_if.wdata1_r\[4\] io_in[4] u_cpu.rf_ram_if.wdata1_r\[3\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06326__A1 _02512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09609_ _00063_ io_in[4] u_cpu.rf_ram.memory\[20\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10881_ _01310_ io_in[4] u_cpu.rf_ram.memory\[25\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06877__A2 _03002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04888__A1 u_cpu.cpu.immdec.imm24_20\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07826__A1 _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06629__A2 _02864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09613__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08251__A1 _03767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10315_ _00748_ io_in[4] u_cpu.rf_ram.memory\[34\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06801__A2 _02955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05396__B _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07167__I _02501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10246_ _00679_ io_in[4] u_cpu.rf_ram.memory\[38\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09763__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06014__B1 u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08554__A2 _04094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10177_ _00623_ io_in[4] u_cpu.rf_ram.memory\[22\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06565__A1 _02748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10740__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08306__A2 _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09503__A1 _04482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06868__A2 _02992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04879__A1 _01402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10890__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06270_ _02512_ _02641_ _02648_ _00104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08490__A1 _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07293__A2 _03235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05150__I _01548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10120__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05221_ _01705_ _01707_ _01709_ _01711_ _01426_ _01712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_129_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08617__I0 u_arbiter.i_wb_cpu_dbus_adr\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05152_ _01398_ _01643_ _01644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06182__S _02578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08242__A1 _03741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07045__A2 _03091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08793__A2 _04227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09960_ _00414_ io_in[4] u_cpu.rf_ram.memory\[54\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05083_ u_cpu.rf_ram.memory\[20\]\[0\] u_cpu.rf_ram.memory\[21\]\[0\] u_cpu.rf_ram.memory\[22\]\[0\]
+ u_cpu.rf_ram.memory\[23\]\[0\] _01572_ _01574_ _01575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_131_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10270__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05151__S1 _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08911_ u_cpu.rf_ram.memory\[96\]\[4\] _04309_ _04314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06910__S _03021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09891_ _00345_ io_in[4] u_cpu.rf_ram.memory\[61\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08842_ _03539_ _04271_ _04272_ _01053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05359__A2 _01848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08773_ _04221_ _01035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05985_ _02305_ _02448_ _02449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07724_ u_cpu.rf_ram.memory\[90\]\[6\] _03475_ _03482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04936_ u_cpu.cpu.ctrl.o_ibus_adr\[5\] _01451_ u_cpu.cpu.ctrl.o_ibus_adr\[6\] _01454_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_38_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07655_ u_cpu.rf_ram.memory\[36\]\[0\] _03442_ _03443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06859__A2 _02992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_04867_ u_cpu.cpu.genblk3.csr.o_new_irq u_cpu.cpu.state.genblk1.misalign_trap_sync_r
+ _01392_ _01393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_92_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06606_ _02752_ _02844_ _02851_ _00237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07586_ _03347_ _03402_ _03404_ _00664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09325_ _04545_ _04546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07808__A1 _03349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06537_ u_cpu.rf_ram.memory\[40\]\[0\] _02812_ _02813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09256_ u_cpu.rf_ram.memory\[85\]\[1\] _04506_ _04508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09636__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08481__A1 _03747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06468_ _01435_ _02765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__08572__S _02445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07284__A2 _03225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05295__A1 _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08207_ u_cpu.cpu.decode.opcode\[1\] _03798_ _03806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05419_ _01597_ _01907_ _01908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09187_ u_cpu.rf_ram.memory\[69\]\[6\] _04459_ _04466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06399_ _02502_ _02718_ _02723_ _00158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10613__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08138_ u_cpu.rf_ram.memory\[113\]\[7\] _03731_ _03739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08233__A1 _03767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07036__A2 _03091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05047__A1 _01419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08784__A2 _04227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09786__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08069_ u_arbiter.i_wb_cpu_dbus_dat\[14\] _03683_ _03696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05142__S1 _01616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10100_ _00546_ io_in[4] u_cpu.rf_ram.memory\[137\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11080_ _11080_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__10763__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08536__A2 _04084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10031_ _00477_ io_in[4] u_cpu.rf_ram.memory\[13\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10933_ _01361_ io_in[4] u_cpu.cpu.state.ibus_cyc vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10864_ _01293_ io_in[4] u_cpu.rf_ram.memory\[27\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10143__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10795_ _01224_ io_in[4] u_cpu.rf_ram.memory\[10\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08472__A1 u_cpu.cpu.immdec.imm19_12_20\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07275__A2 _03225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05286__A1 _01399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[56\] u_scanchain_local.module_data_in\[55\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[18\] u_scanchain_local.clk u_scanchain_local.module_data_in\[56\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_144_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10293__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08224__A1 _03791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07027__A2 _03081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05133__S1 _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06786__A1 _02752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10229_ _00019_ io_in[4] u_cpu.rf_ram_if.rdata1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06538__A1 _02738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05573__C _01426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05770_ u_cpu.rf_ram.memory\[108\]\[7\] u_cpu.rf_ram.memory\[109\]\[7\] u_cpu.rf_ram.memory\[110\]\[7\]
+ u_cpu.rf_ram.memory\[111\]\[7\] _01598_ _01573_ _02255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_47_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07440_ u_cpu.rf_ram.memory\[131\]\[4\] _03315_ _03320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09659__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05513__A2 _02000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06710__A1 _02748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07371_ _03169_ _03275_ _03281_ _00572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09110_ _04288_ _04419_ _04423_ _01170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10636__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06322_ _02502_ _02673_ _02678_ _00126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08463__A1 _03825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05277__A1 _01636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09041_ u_cpu.rf_ram.memory\[104\]\[5\] _04379_ _04385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06253_ _02468_ _02637_ _02638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_136_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05204_ u_cpu.rf_ram.memory\[8\]\[1\] u_cpu.rf_ram.memory\[9\]\[1\] u_cpu.rf_ram.memory\[10\]\[1\]
+ u_cpu.rf_ram.memory\[11\]\[1\] _01546_ _01550_ _01695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_129_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08215__A1 _03773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07018__A2 _03081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06184_ u_cpu.rf_ram_if.wdata0_r\[6\] u_cpu.rf_ram_if.wdata1_r\[6\] _02478_ _02595_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05029__A1 _01445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10786__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05135_ _01541_ _01625_ _01626_ _01627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_144_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05066_ u_cpu.rf_ram.memory\[12\]\[0\] u_cpu.rf_ram.memory\[13\]\[0\] u_cpu.rf_ram.memory\[14\]\[0\]
+ u_cpu.rf_ram.memory\[15\]\[0\] _01556_ _01557_ _01558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09943_ _00397_ io_in[4] u_cpu.rf_ram.memory\[56\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08518__A2 _03988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10016__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09874_ _00328_ io_in[4] u_cpu.rf_ram.memory\[63\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06529__A1 _02750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08825_ _04237_ _04254_ _04258_ _01050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08756_ _04212_ _01027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05968_ u_cpu.cpu.state.init_done _02433_ _02434_ _02435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_72_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07471__S _03334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10166__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07707_ _03357_ _03465_ _03472_ _00717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_04919_ _01429_ u_cpu.cpu.state.ibus_cyc _01441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08687_ _04172_ _00998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_05899_ _02379_ _02380_ _02381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07638_ _03343_ _03432_ _03433_ _00687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07569_ u_cpu.rf_ram.memory\[125\]\[2\] _03392_ _03395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09308_ u_cpu.rf_ram.memory\[111\]\[0\] _04536_ _04537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10580_ _01010_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05268__A1 _01553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05807__A3 _02291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09239_ _04498_ _01224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08206__A1 _03761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07009__A2 _03071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06768__A1 _02752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05440__A1 _01645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08509__A2 _03668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11063_ _11063_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__05674__B _01416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05991__A2 u_cpu.cpu.immdec.imm11_7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10014_ _00460_ io_in[4] u_cpu.rf_ram.memory\[141\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09182__A2 _04459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10509__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[1\] u_cpu.cpu.genblk3.csr.i_mtip io_in[3] u_arbiter.o_wb_cpu_we
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_ack vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_95_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06940__A1 _02684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09801__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10659__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10916_ _01345_ io_in[4] u_cpu.rf_ram.memory\[89\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07496__A2 _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10847_ _01276_ io_in[4] u_cpu.rf_ram.memory\[88\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09951__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08445__A1 _01373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07248__A2 _03206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10778_ _01207_ io_in[4] u_cpu.rf_ram.memory\[84\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08996__A2 _04359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10039__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08748__A2 _02682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06460__S _02756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07420__A2 _03305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06940_ _02684_ _02695_ _03040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10189__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09173__A2 _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06871_ u_cpu.rf_ram.memory\[60\]\[0\] _03002_ _03003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07184__A1 _03161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05822_ u_arbiter.i_wb_cpu_dbus_we _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08610_ _04127_ _00966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09590_ _00044_ io_in[4] u_cpu.rf_ram.memory\[81\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06931__A1 _02961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08541_ _03553_ _04084_ _04091_ _00933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_u_scanchain_local.scan_flop\[4\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05753_ _01540_ _02237_ _01564_ _02238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_36_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08472_ u_cpu.cpu.immdec.imm19_12_20\[5\] _03798_ _04016_ _04036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05684_ u_cpu.rf_ram.memory\[104\]\[6\] u_cpu.rf_ram.memory\[105\]\[6\] u_cpu.rf_ram.memory\[106\]\[6\]
+ u_cpu.rf_ram.memory\[107\]\[6\] _01615_ _01616_ _02170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_35_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07487__A2 _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08684__B2 u_cpu.cpu.ctrl.o_ibus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05498__A1 _01397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07423_ _03167_ _03305_ _03310_ _00595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07354_ u_cpu.rf_ram.memory\[136\]\[6\] _03265_ _03272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08436__A1 _03744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07239__A2 _03206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08436__B2 _03778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09484__I0 _02596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06305_ _02507_ _02662_ _02668_ _00119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08987__A2 _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07285_ _03173_ _03225_ _03233_ _00534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05345__S1 _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09024_ _04292_ _04369_ _04375_ _01132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06236_ u_cpu.rf_ram.memory\[78\]\[0\] _02628_ _02629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09236__I0 _02573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08739__A2 _04199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06167_ _02582_ _00067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05118_ _01544_ _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07411__A2 _03295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06098_ _02464_ _02521_ _02539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05049_ _01540_ _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09926_ _00380_ io_in[4] u_cpu.rf_ram.memory\[58\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09164__A2 _04449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09824__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09857_ _00311_ io_in[4] u_cpu.rf_ram.memory\[64\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07175__A1 _03171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08911__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08808_ _03761_ _03778_ _03779_ _03788_ _04243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_73_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09788_ _00242_ io_in[4] u_cpu.rf_ram.memory\[77\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06922__A1 _02638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10801__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05281__S0 _01680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08739_ _03547_ _04199_ _04203_ _01019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09974__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05489__A1 _01594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10701_ _01130_ io_in[4] u_cpu.rf_ram.memory\[103\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10951__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06150__A2 _02563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10632_ _01061_ io_in[4] u_cpu.rf_ram.memory\[94\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08978__A2 _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10563_ _00993_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05669__B _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05336__S1 _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06989__A1 _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10494_ _00927_ io_in[4] u_cpu.rf_ram.memory\[32\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07650__A2 _03432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05388__C _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07402__A2 _03295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10331__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_scanchain_local.scan_flop\[19\] u_arbiter.i_wb_cpu_rdt\[16\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[13\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_49_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11046_ _11046_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__09155__A2 _04197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07166__A1 _03165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08363__C2 _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10481__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05272__S0 _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06141__A2 _02563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08418__A1 _03802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07070_ _02584_ u_cpu.rf_ram.memory\[15\]\[2\] _03109_ _03112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07641__A2 _03432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06021_ u_cpu.rf_ram_if.genblk1.wtrig0_r _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09847__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06190__S _02578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[52\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06452__I0 _02573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07972_ _03539_ _03626_ _03627_ _00828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10824__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09711_ _00165_ io_in[4] u_cpu.rf_ram.memory\[47\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09146__A2 _04439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06923_ _03030_ _03031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07157__A1 _03157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09997__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09642_ _00096_ io_in[4] u_cpu.rf_ram.memory\[78\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06854_ _02953_ _02992_ _02993_ _00343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06904__A1 _02969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[67\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05263__S0 _01646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05805_ _01553_ _02289_ _01648_ _02290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09573_ _00027_ io_in[4] u_cpu.rf_ram.memory\[82\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06785_ u_cpu.rf_ram.memory\[64\]\[6\] _02944_ _02951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08106__B1 _03718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06380__A2 _02708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08524_ u_cpu.cpu.genblk3.csr.mie_mtie u_cpu.cpu.genblk3.csr.mstatus_mie u_cpu.cpu.genblk3.csr.i_mtip
+ _04081_ _04082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_05736_ u_cpu.rf_ram.memory\[4\]\[7\] u_cpu.rf_ram.memory\[5\]\[7\] u_cpu.rf_ram.memory\[6\]\[7\]
+ u_cpu.rf_ram.memory\[7\]\[7\] _01578_ _01580_ _02221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_36_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08455_ u_cpu.cpu.immdec.imm19_12_20\[3\] _03797_ _04015_ _04021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05667_ _01636_ _02152_ _02153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06132__A2 _02551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10204__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07406_ u_cpu.rf_ram.memory\[133\]\[5\] _03295_ _03301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08386_ _03761_ _03860_ _03941_ _03959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08409__A1 _03776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07880__A2 _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05598_ u_cpu.rf_ram.memory\[100\]\[5\] u_cpu.rf_ram.memory\[101\]\[5\] u_cpu.rf_ram.memory\[102\]\[5\]
+ u_cpu.rf_ram.memory\[103\]\[5\] _01577_ _01549_ _02085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_11_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05891__A1 _02361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07337_ _03171_ _03255_ _03262_ _00557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09082__A1 _04296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05489__B _01564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08580__S _02445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07268_ _02638_ _02832_ _03224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07632__A2 _03422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10354__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05643__A1 _01406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06219_ _02492_ _02614_ _02617_ _00084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09007_ u_cpu.rf_ram.memory\[102\]\[6\] _04359_ _04366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06691__I0 _02590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07199_ u_cpu.rf_ram.memory\[71\]\[0\] _03186_ _03187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09137__A2 _02682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09909_ _00363_ io_in[4] u_cpu.rf_ram.memory\[19\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07699__A2 _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08896__A1 _04292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08648__A1 u_cpu.rf_ram.memory\[30\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08755__S _04208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06123__A2 _02551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07871__A2 _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05882__A1 _01369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10615_ _01044_ io_in[4] u_cpu.rf_ram.memory\[93\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07623__A2 _03422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08820__A1 u_cpu.cpu.immdec.imm11_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10546_ _00978_ io_in[4] u_cpu.rf_ram.memory\[30\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05634__A1 _01399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10477_ _00910_ io_in[4] u_cpu.cpu.immdec.imm30_25\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10847__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07387__A1 _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09128__A2 _04429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11029_ _11029_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_110_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05165__A3 _01656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06362__A2 _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10227__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06570_ u_cpu.rf_ram.memory\[119\]\[7\] _02823_ _02831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08639__A1 _03539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05153__I _01540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05521_ u_cpu.rf_ram.memory\[116\]\[4\] u_cpu.rf_ram.memory\[117\]\[4\] u_cpu.rf_ram.memory\[118\]\[4\]
+ u_cpu.rf_ram.memory\[119\]\[4\] _01623_ _01624_ _02009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_61_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09300__A2 _04526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06114__A2 _02541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07311__A1 _03163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08240_ _02333_ _03740_ _03834_ _00889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05452_ u_cpu.rf_ram.memory\[76\]\[3\] u_cpu.rf_ram.memory\[77\]\[3\] u_cpu.rf_ram.memory\[78\]\[3\]
+ u_cpu.rf_ram.memory\[79\]\[3\] _01577_ _01549_ _01941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_60_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07862__A2 _03558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10377__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08171_ _03754_ _03755_ _03770_ _03771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09064__A1 _04296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05383_ _01554_ _01871_ _01417_ _01872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_20_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07122_ u_cpu.rf_ram.memory\[140\]\[1\] _03139_ _03141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07614__A2 _03412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05625__A1 _01553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07053_ _02584_ u_cpu.rf_ram.memory\[9\]\[2\] _03100_ _03103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06004_ u_cpu.cpu.immdec.imm11_7\[1\] _02460_ _02461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05928__A2 _02406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09119__A2 _04197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07955_ u_cpu.rf_ram.memory\[115\]\[1\] _03616_ _03618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08327__B1 _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06906_ _02573_ u_cpu.rf_ram.memory\[5\]\[0\] _03021_ _03022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07886_ _02584_ u_cpu.rf_ram.memory\[8\]\[2\] _03577_ _03580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09625_ _00079_ io_in[4] u_cpu.rf_ram.memory\[7\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06837_ u_cpu.rf_ram.memory\[62\]\[1\] _02982_ _02984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07550__A1 _03347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06353__A2 _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09556_ u_cpu.rf_ram.memory\[23\]\[6\] _04674_ _04681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05063__I _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06768_ _02752_ _02934_ _02941_ _00309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_70_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08507_ _03741_ _03988_ _04067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05719_ _01539_ _02195_ _02204_ _02205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_23_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06105__A2 _02541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09487_ _04642_ _01328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06699_ _02561_ _02626_ _02903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08438_ _03754_ _04002_ _04006_ _04007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07853__A2 _03558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08369_ _03773_ _03858_ _03942_ _03943_ _03944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_7_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10400_ _00833_ io_in[4] u_cpu.rf_ram.memory\[116\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07605__A2 _03412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05616__A1 _01645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10331_ _00764_ io_in[4] u_cpu.rf_ram.memory\[120\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09358__A2 _04556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10262_ _00695_ io_in[4] u_cpu.rf_ram.memory\[36\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07369__A1 _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10193_ _00639_ io_in[4] u_cpu.rf_ram.memory\[127\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05919__A2 _02313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06041__A1 _02460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09530__A2 _04664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06344__A2 _02686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08097__A2 _03653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07844__A2 _03541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09692__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05855__A1 u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09046__A1 _04296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10529_ _00962_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09349__A2 _04556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06280__A1 _02492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07080__I0 _02599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07780__A1 _03357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06583__A2 _02834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04952_ u_cpu.cpu.ctrl.o_ibus_adr\[9\] _01464_ _01467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07740_ _02333_ _03494_ _03495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_111_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07907__I0 _02590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09521__A2 _04654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04883_ _01370_ u_cpu.cpu.bne_or_bge _01409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07671_ _02311_ _02773_ _03451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07532__A1 _03347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05138__A3 _01629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06335__A2 _02686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09410_ _04478_ _04595_ _04600_ _01293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06622_ _02750_ _02854_ _02860_ _00244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_19_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06908__S _03021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09341_ _04484_ _04546_ _04554_ _01270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__04897__A2 _01368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06553_ _02473_ _02683_ _02821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09285__A1 _04482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08088__A2 _03683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06099__A1 _02475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05504_ _01422_ _01982_ _01991_ _01992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_09272_ u_cpu.rf_ram.memory\[110\]\[0\] _04516_ _04517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06484_ _01408_ _01370_ _02779_ _02780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__07835__A2 _03541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05846__A1 _02305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05435_ _01917_ _01919_ _01921_ _01923_ _01607_ _01924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_08223_ _03818_ _03819_ _03790_ _03810_ _03820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_119_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08154_ _02765_ u_arbiter.i_wb_cpu_rdt\[0\] _03753_ _03754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_u_scanchain_local.scan_flop\[20\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05366_ _01849_ _01851_ _01853_ _01855_ _01568_ _01856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__07599__A1 _02706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07105_ _02957_ _03129_ _03131_ _00456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08085_ u_arbiter.i_wb_cpu_dbus_dat\[20\] _03683_ _03706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08260__A2 _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05297_ _01554_ _01786_ _01787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07036_ u_cpu.rf_ram.memory\[52\]\[2\] _03091_ _03094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06442__I _02506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08012__A2 _01442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05058__I _01549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05457__S0 _01680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08987_ u_cpu.rf_ram.memory\[101\]\[5\] _04349_ _04355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07938_ _03543_ _03606_ _03608_ _00813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09512__A2 _04654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10542__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07869_ u_cpu.rf_ram.memory\[121\]\[2\] _03568_ _03571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06326__A2 _02673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08720__B1 _04175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09608_ _00062_ io_in[4] u_cpu.rf_ram.memory\[20\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10880_ _01309_ io_in[4] u_cpu.rf_ram.memory\[25\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__04888__A2 _01387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09539_ _04482_ _04664_ _04671_ _01351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10692__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07826__A2 _03541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09028__A1 _04296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08251__A2 _03774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06262__A1 _02492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10314_ _00747_ io_in[4] u_cpu.rf_ram.memory\[35\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_4_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09908__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08003__A2 _03636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10245_ _00014_ io_in[4] u_cpu.rf_ram_if.rdata0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10072__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06014__A1 u_cpu.rf_ram_if.genblk1.wtrig0_r vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05448__S0 _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10176_ _00622_ io_in[4] u_cpu.rf_ram.memory\[12\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06565__A2 _02823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07762__A1 _03357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09503__A2 _04644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06317__A2 _02673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07514__A1 _03347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04879__A2 _01404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09267__A1 _04482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07817__A2 _03530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[43\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08943__S _04331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05220_ _01542_ _01710_ _01418_ _01711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05151_ u_cpu.rf_ram.memory\[124\]\[0\] u_cpu.rf_ram.memory\[125\]\[0\] u_cpu.rf_ram.memory\[126\]\[0\]
+ u_cpu.rf_ram.memory\[127\]\[0\] _01545_ _01642_ _01643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_7_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08242__A2 _03818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10415__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05082_ _01573_ _01574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09588__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08910_ _04288_ _04309_ _04313_ _01080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09890_ _00344_ io_in[4] u_cpu.rf_ram.memory\[61\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06005__A1 _02460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05439__S0 _01646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07053__I0 _02584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08841_ u_cpu.rf_ram.memory\[97\]\[0\] _04271_ _04272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10565__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06556__A2 _02823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07753__A1 u_cpu.rf_ram.memory\[92\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08772_ _02587_ u_cpu.rf_ram.memory\[2\]\[3\] _04217_ _04221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05984_ _02447_ _02365_ _02448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07723_ _03355_ _03475_ _03481_ _00724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04935_ _01445_ _01452_ _01453_ u_arbiter.o_wb_cpu_adr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06308__A2 _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07505__A1 _03357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08702__B1 _04175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07654_ _03441_ _03442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_04866_ _01378_ _01383_ _01392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_81_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06605_ u_cpu.rf_ram.memory\[139\]\[6\] _02844_ _02851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07585_ u_cpu.rf_ram.memory\[124\]\[1\] _03402_ _03404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09324_ _02475_ _02602_ _04545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06536_ _02811_ _02812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07808__A2 _03530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05819__A1 _01406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09255_ _04468_ _04506_ _04507_ _01231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06467_ _02764_ _00185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08481__A2 _03825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07469__S _03334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05295__A2 _01784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08206_ _03761_ _03782_ _03804_ _03805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06492__A1 _01680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05418_ u_cpu.rf_ram.memory\[108\]\[3\] u_cpu.rf_ram.memory\[109\]\[3\] u_cpu.rf_ram.memory\[110\]\[3\]
+ u_cpu.rf_ram.memory\[111\]\[3\] _01598_ _01573_ _01907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_06398_ u_cpu.rf_ram.memory\[48\]\[4\] _02718_ _02723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09186_ _04292_ _04459_ _04465_ _01204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08137_ _03553_ _03731_ _03738_ _00882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05349_ u_cpu.rf_ram.memory\[92\]\[2\] u_cpu.rf_ram.memory\[93\]\[2\] u_cpu.rf_ram.memory\[94\]\[2\]
+ u_cpu.rf_ram.memory\[95\]\[2\] _01610_ _01611_ _01839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10095__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09430__A1 _04480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08233__A2 _03778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05047__A2 _01420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08068_ _03694_ _03695_ _00856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07992__A1 _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10908__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06795__A2 _02955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07019_ _02959_ _03081_ _03084_ _00417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10030_ _00476_ io_in[4] u_cpu.rf_ram.memory\[13\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06547__A2 _02812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09497__A1 _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10932_ _01360_ io_in[4] u_cpu.rf_ram.memory\[23\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[66\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10863_ _01292_ io_in[4] u_cpu.rf_ram.memory\[27\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08763__S _04208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10794_ _01223_ io_in[4] u_cpu.rf_ram.memory\[10\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08472__A2 _03798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10438__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09730__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[49\] u_scanchain_local.module_data_in\[48\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[11\] u_scanchain_local.clk u_scanchain_local.module_data_in\[49\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_67_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05200__B _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10588__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06786__A2 _02944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09880__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10228_ _00018_ io_in[4] u_cpu.rf_ram_if.rdata1\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06538__A2 _02812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10159_ _00605_ io_in[4] u_cpu.rf_ram.memory\[131\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09488__A1 _02469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05870__B _01369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05349__I0 u_cpu.rf_ram.memory\[92\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06458__S _02756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08160__A1 _01435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06710__A2 _02904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07370_ u_cpu.rf_ram.memory\[135\]\[5\] _03275_ _03281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06321_ u_cpu.rf_ram.memory\[44\]\[4\] _02673_ _02678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08463__A2 _03776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09040_ _04290_ _04379_ _04384_ _01139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06474__A1 _02311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06252_ _02459_ _02623_ _02637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05203_ _01406_ _01631_ _01694_ _00000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06183_ _02594_ _00071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_11_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09412__A1 _04480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08215__A2 _03810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05134_ _01564_ _01626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07974__A1 _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06777__A2 _02944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09942_ _00396_ io_in[4] u_cpu.rf_ram.memory\[56\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05065_ _01548_ _01557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09873_ _00327_ io_in[4] u_cpu.rf_ram.memory\[63\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06529__A2 _02801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08774__I0 _02590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08824_ u_cpu.cpu.immdec.imm11_7\[2\] _04237_ _04257_ _03740_ _04258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_58_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08755_ _02587_ u_cpu.rf_ram.memory\[3\]\[3\] _04208_ _04212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_85_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05967_ _01372_ _01374_ _02434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07706_ u_cpu.rf_ram.memory\[91\]\[6\] _03465_ _03472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04918_ _01431_ _01439_ _01440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08686_ u_cpu.cpu.ctrl.o_ibus_adr\[14\] _04155_ _04157_ u_cpu.cpu.ctrl.o_ibus_adr\[15\]
+ _04172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_26_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09603__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08151__A1 _02765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05898_ u_arbiter.i_wb_cpu_ibus_adr\[0\] u_cpu.cpu.ctrl.pc_plus_4_cy_r _02380_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07637_ u_cpu.rf_ram.memory\[37\]\[0\] _03432_ _03433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04849_ _01374_ _01375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_53_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05504__A3 _01991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06701__A2 _02904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07568_ _03347_ _03392_ _03394_ _00656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09307_ _04535_ _04536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06519_ _02738_ _02801_ _02802_ _00199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09753__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07499_ _03353_ _03345_ _03354_ _00627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05268__A2 _01758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09238_ _02581_ u_cpu.rf_ram.memory\[10\]\[1\] _04496_ _04498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10730__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09169_ u_cpu.rf_ram.memory\[108\]\[6\] _04449_ _04456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08206__A2 _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06217__A1 _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06768__A2 _02934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10880__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05440__A2 _01928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11062_ _11062_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_7_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07717__A1 _03349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05991__A3 u_cpu.cpu.immdec.imm11_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10013_ _00459_ io_in[4] u_cpu.rf_ram.memory\[141\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07193__A2 _03176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10110__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06940__A2 _02695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__04951__A1 _01445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10915_ _01344_ io_in[4] u_cpu.rf_ram.memory\[100\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10260__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10846_ _01275_ io_in[4] u_cpu.rf_ram.memory\[88\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10777_ _01206_ io_in[4] u_cpu.rf_ram.memory\[69\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08445__A2 u_cpu.cpu.decode.opcode\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08225__C _03797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07256__I0 _02584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07956__A1 _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06759__A2 _02934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05982__A3 _02401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06870_ _03001_ _03002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09626__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05156__I _01416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07184__A2 _03176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05821_ _02304_ _02305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06931__A2 _03031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08540_ u_cpu.rf_ram.memory\[32\]\[6\] _04084_ _04091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06188__S _02460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05752_ u_cpu.rf_ram.memory\[48\]\[7\] u_cpu.rf_ram.memory\[49\]\[7\] u_cpu.rf_ram.memory\[50\]\[7\]
+ u_cpu.rf_ram.memory\[51\]\[7\] _01544_ _01548_ _02237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_78_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10603__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08133__A1 _03549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08471_ _03768_ _03774_ _04034_ _03740_ _04035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05683_ _01597_ _02168_ _02169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09776__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08684__A2 _04155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05498__A2 _01985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07422_ u_cpu.rf_ram.memory\[132\]\[4\] _03305_ _03310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06916__S _03021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10753__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07353_ _03169_ _03265_ _03271_ _00564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08436__A2 _03818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08416__B _03741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06304_ u_cpu.rf_ram.memory\[45\]\[5\] _02662_ _02668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06447__A1 _02752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07284_ u_cpu.rf_ram.memory\[138\]\[7\] _03225_ _03233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06998__A2 _03071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09023_ u_cpu.rf_ram.memory\[103\]\[5\] _04369_ _04375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06235_ _02627_ _02628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_129_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05670__A2 _02151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06166_ _02581_ u_cpu.rf_ram.memory\[1\]\[1\] _02578_ _02582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_102_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05117_ _01540_ _01609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06097_ _02517_ _02530_ _02538_ _00041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05048_ _01389_ _01391_ _01395_ _01540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_09925_ _00379_ io_in[4] u_cpu.rf_ram.memory\[58\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10133__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05494__C _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09856_ _00310_ io_in[4] u_cpu.rf_ram.memory\[65\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08578__S _02445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07175__A2 _03159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08372__A1 _02436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08807_ _03747_ _03825_ _04000_ _04241_ _03782_ _04242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_58_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05186__A1 _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09787_ _00241_ io_in[4] u_cpu.rf_ram.memory\[77\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06999_ _02957_ _03071_ _03073_ _00408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06922__A2 _02684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10283__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08738_ u_cpu.rf_ram.memory\[109\]\[3\] _04199_ _04203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05281__S1 _01681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08669_ _04163_ _00989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_26_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10700_ _01129_ io_in[4] u_cpu.rf_ram.memory\[103\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05489__A2 _01976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10631_ _01060_ io_in[4] u_cpu.rf_ram.memory\[97\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08427__A2 _02438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08326__B _03906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06438__A1 _02746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10562_ _00992_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06989__A2 _03061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10493_ _00926_ io_in[4] u_cpu.cpu.genblk3.csr.timer_irq_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05661__A2 _02142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07938__A1 _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05685__B _01416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09649__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11114_ u_scanchain_local.data_out io_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11045_ _11045_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_122_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08488__S _01436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10626__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08363__A1 u_cpu.cpu.immdec.imm24_20\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07166__A2 _03159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08363__B2 u_cpu.cpu.immdec.imm30_25\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09799__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.output_buffers\[3\]_I u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05272__S1 _01652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08115__A1 u_arbiter.i_wb_cpu_rdt\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10776__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08666__A2 _04155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10829_ _01258_ io_in[4] u_cpu.rf_ram.memory\[111\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08418__A2 _03826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10006__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06429__A1 _02738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07477__I0 _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08951__S _04331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09091__A2 _04409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05101__A1 _01589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09993__D _00000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06020_ _02476_ _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10156__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07971_ u_cpu.rf_ram.memory\[116\]\[0\] _03626_ _03627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09710_ _00164_ io_in[4] u_cpu.rf_ram.memory\[47\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06922_ _02638_ _02684_ _03030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08354__A1 _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07157__A2 _03159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09641_ _00095_ io_in[4] u_cpu.rf_ram.memory\[78\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06853_ u_cpu.rf_ram.memory\[61\]\[0\] _02992_ _02993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06904__A2 _03012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05804_ u_cpu.rf_ram.memory\[76\]\[7\] u_cpu.rf_ram.memory\[77\]\[7\] u_cpu.rf_ram.memory\[78\]\[7\]
+ u_cpu.rf_ram.memory\[79\]\[7\] _01577_ _01549_ _02289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_55_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05263__S1 _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09572_ _00026_ io_in[4] u_cpu.rf_ram.memory\[82\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06784_ _02750_ _02944_ _02950_ _00316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08106__A1 u_arbiter.i_wb_cpu_rdt\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08523_ _02311_ _02448_ _04081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_64_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05735_ _01398_ _02219_ _01417_ _02220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_91_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06668__A1 _02742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08454_ u_cpu.cpu.immdec.imm19_12_20\[2\] _04020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05666_ u_cpu.rf_ram.memory\[60\]\[6\] u_cpu.rf_ram.memory\[61\]\[6\] u_cpu.rf_ram.memory\[62\]\[6\]
+ u_cpu.rf_ram.memory\[63\]\[6\] _01598_ _01573_ _02152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_17_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07405_ _03167_ _03295_ _03300_ _00587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05340__A1 _01398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08385_ _03858_ _03943_ _03958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08409__A2 _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05597_ _01594_ _02083_ _01416_ _02084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06445__I _02511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05891__A2 _02372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07336_ u_cpu.rf_ram.memory\[49\]\[6\] _03255_ _03262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09082__A2 _04399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07093__A1 _02963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07267_ _03223_ _00526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09006_ _04292_ _04359_ _04365_ _01124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07477__S _03334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06218_ u_cpu.rf_ram.memory\[80\]\[2\] _02614_ _02617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06840__A1 _02959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05643__A2 _02080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07198_ _03185_ _03186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_104_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06149_ u_cpu.rf_ram.memory\[20\]\[5\] _02563_ _02569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10649__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07396__A2 _03295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09941__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09908_ _00362_ io_in[4] u_cpu.rf_ram.memory\[19\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_101_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08345__B2 _03877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05159__A1 _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09839_ _00293_ io_in[4] u_cpu.rf_ram.memory\[67\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10799__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08896__A2 _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__04906__A1 _01429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08648__A2 _04145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10029__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07320__A2 _03245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05331__A1 _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10614_ _01043_ io_in[4] u_cpu.rf_ram.memory\[93\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05882__A2 _01370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09073__A2 _04399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10179__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10545_ _00977_ io_in[4] u_cpu.rf_ram.memory\[30\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08820__A2 _03798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05634__A2 _02120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10476_ _00909_ io_in[4] u_cpu.cpu.immdec.imm30_25\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05190__S0 _01680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08959__I0 u_arbiter.i_wb_cpu_rdt\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[31\] u_arbiter.i_wb_cpu_rdt\[28\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[25\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__08503__C _03797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07387__A2 _03285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11028_ _11028_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_77_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08887__A2 _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06898__A1 _02963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05570__A1 _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08639__A2 _04145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05520_ _01541_ _02007_ _02008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06466__S _02756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07311__A2 _03245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05322__A1 _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05451_ _01667_ _01939_ _01940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08170_ _03765_ _03769_ _03770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09814__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05382_ u_cpu.rf_ram.memory\[12\]\[3\] u_cpu.rf_ram.memory\[13\]\[3\] u_cpu.rf_ram.memory\[14\]\[3\]
+ u_cpu.rf_ram.memory\[15\]\[3\] _01556_ _01557_ _01871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09064__A2 _04389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07121_ _02953_ _03139_ _03140_ _00463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07052_ _03102_ _00432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06822__A1 _02959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05181__S0 _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06003_ u_cpu.rf_ram_if.genblk1.wtrig0_r _02460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_12_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09964__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07378__A2 _03285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10941__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06050__A2 _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07954_ _03539_ _03616_ _03617_ _00820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08327__A1 _03763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08327__B2 _03744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07824__I _02486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06905_ _02524_ _02577_ _03021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07885_ _03579_ _00789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08878__A2 _04282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09624_ _00078_ io_in[4] u_cpu.rf_ram.memory\[7\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06836_ _02953_ _02982_ _02983_ _00335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07550__A2 _03382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09555_ _04480_ _04674_ _04680_ _01358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05561__A1 _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06767_ u_cpu.rf_ram.memory\[65\]\[6\] _02934_ _02941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08506_ _04016_ _04064_ _04065_ _04066_ _00923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_05718_ _02197_ _02199_ _02201_ _02203_ _01568_ _02204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_19_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09486_ _02599_ u_cpu.rf_ram.memory\[0\]\[7\] _04634_ _04642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06698_ _02902_ _00278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07302__A2 _03235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10321__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08437_ _03999_ _03988_ _04003_ _04005_ _03801_ _04006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_106_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05649_ _01554_ _02134_ _02135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05313__A1 _01594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05864__A2 _02324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08368_ _03831_ _03861_ _03902_ _03943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08591__S _04115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09055__A2 _04389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07319_ _03171_ _03245_ _03252_ _00549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08299_ u_cpu.rf_ram.memory\[114\]\[4\] _03879_ _03884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08802__A2 _03797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10471__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05616__A2 _02102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10330_ _00763_ io_in[4] u_cpu.rf_ram.memory\[117\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05172__S0 _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08015__B1 _03654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10261_ _00694_ io_in[4] u_cpu.rf_ram.memory\[37\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07369__A2 _03275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10192_ _00638_ io_in[4] u_cpu.rf_ram.memory\[128\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08869__A2 _04282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08766__S _04217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07541__A2 _03372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05552__A1 _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09837__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09294__A2 _04526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05304__A1 _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[51\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10814__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09046__A2 _04379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09987__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06804__A1 u_cpu.rf_ram.memory\[29\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10528_ _00961_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_u_scanchain_local.scan_flop\[66\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06280__A2 _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10459_ _00892_ io_in[4] u_cpu.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08557__A1 _03551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06032__A2 _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07780__A2 _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04951_ _01445_ _01465_ _01466_ u_arbiter.o_wb_cpu_adr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07670_ _03359_ _03442_ _03450_ _00702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_93_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04882_ _01369_ _01408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_93_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07532__A2 _03372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10344__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06621_ u_cpu.rf_ram.memory\[77\]\[5\] _02854_ _02860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05543__A1 _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09340_ u_cpu.rf_ram.memory\[87\]\[7\] _04546_ _04554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06552_ _02754_ _02812_ _02820_ _00214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09285__A2 _04516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05503_ _01984_ _01986_ _01988_ _01990_ _01628_ _01991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_61_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09271_ _04515_ _04516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06099__A2 _02539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[19\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06483_ _02771_ _02778_ _02779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10494__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08222_ _03741_ _03742_ _03819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05434_ _01614_ _01922_ _01654_ _01923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_14_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09037__A2 _04379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07048__A1 _02577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08245__B1 _03801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08153_ _01436_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[0\] _03753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_20_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05365_ _01636_ _01854_ _01417_ _01855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_101_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08424__B u_cpu.cpu.decode.opcode\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07599__A2 _02821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07104_ u_cpu.rf_ram.memory\[141\]\[1\] _03129_ _03131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07819__I _02481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08084_ _03704_ _03705_ _00862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05767__C _01628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05296_ u_cpu.rf_ram.memory\[4\]\[2\] u_cpu.rf_ram.memory\[5\]\[2\] u_cpu.rf_ram.memory\[6\]\[2\]
+ u_cpu.rf_ram.memory\[7\]\[2\] _01546_ _01550_ _01786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_49_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07035_ _02957_ _03091_ _03093_ _00424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06271__A2 _02641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06023__A2 _02460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07220__A1 _03161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05457__S1 _01681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08986_ _04290_ _04349_ _04354_ _01115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07771__A2 _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07937_ u_cpu.rf_ram.memory\[122\]\[1\] _03606_ _03608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05782__A1 _01601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07868_ _03543_ _03568_ _03570_ _00781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07523__A2 _03362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06819_ u_cpu.rf_ram.memory\[63\]\[1\] _02972_ _02974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09607_ _00061_ io_in[4] u_cpu.rf_ram.memory\[20\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07799_ u_cpu.rf_ram.memory\[34\]\[7\] _03520_ _03528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09538_ u_cpu.rf_ram.memory\[89\]\[6\] _04664_ _04671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10837__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09276__A2 _04516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09469_ u_cpu.rf_ram.memory\[24\]\[7\] _04625_ _04633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09028__A2 _04369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05393__S0 _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07039__A1 _02961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08787__A1 _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08334__B _02305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05145__S0 _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10313_ _00746_ io_in[4] u_cpu.rf_ram.memory\[35\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06262__A2 _02641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10217__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[4\]_D u_arbiter.i_wb_cpu_rdt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08539__A1 _03551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10244_ _00013_ io_in[4] u_cpu.rf_ram_if.rdata0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09200__A2 _04470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05448__S1 _01652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10175_ _00621_ io_in[4] u_cpu.rf_ram.memory\[12\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07762__A2 _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10367__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05773__A1 _01594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07514__A2 _03362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09267__A2 _04506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09019__A2 _04369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05384__S0 _01546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08244__B _03835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05150_ _01548_ _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05081_ _01548_ _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08840_ _04270_ _04271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10940__D u_cpu.cpu.o_wdata0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06005__A2 _01412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07202__A1 _03161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05439__S1 _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07753__A2 _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08771_ _04220_ _01034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05764__A1 _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05983_ u_cpu.cpu.genblk3.csr.o_new_irq u_cpu.cpu.state.init_done _02447_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07722_ u_cpu.rf_ram.memory\[90\]\[5\] _03475_ _03481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_04934_ u_arbiter.i_wb_cpu_dbus_adr\[5\] _01443_ _01453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07505__A2 _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07653_ _02561_ _02639_ _03441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05516__A1 _01398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04865_ _01390_ u_cpu.rf_ram_if.rtrig0 _01391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08419__B _03988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06604_ _02750_ _02844_ _02850_ _00236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07584_ _03343_ _03402_ _03403_ _00663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09258__A2 _04506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09323_ _04484_ _04536_ _04544_ _01262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06535_ _02639_ _02810_ _02811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09254_ u_cpu.rf_ram.memory\[85\]\[0\] _04506_ _04507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06466_ _02599_ u_cpu.rf_ram.memory\[4\]\[7\] _02756_ _02764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__05375__S0 _01687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08205_ _03801_ _03803_ _03804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05417_ _01539_ _01877_ _01886_ _01905_ _01906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_09185_ u_cpu.rf_ram.memory\[69\]\[5\] _04459_ _04465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06397_ _02497_ _02718_ _02722_ _00157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08136_ u_cpu.rf_ram.memory\[113\]\[6\] _03731_ _03738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05348_ _01422_ _01828_ _01837_ _01838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09430__A2 _04605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06244__A2 _02628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07441__A1 _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08067_ u_arbiter.i_wb_cpu_rdt\[12\] _03669_ _03678_ u_arbiter.i_wb_cpu_dbus_dat\[12\]
+ _03695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_88_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05279_ _01539_ _01760_ _01769_ _01770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__07992__A2 _03636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07018_ u_cpu.rf_ram.memory\[53\]\[2\] _03081_ _03084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09682__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08941__A1 _04296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05755__A1 _01636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08969_ u_arbiter.i_wb_cpu_rdt\[29\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[13\]
+ _04331_ _04345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_25_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09497__A2 _04644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10931_ _01359_ io_in[4] u_cpu.rf_ram.memory\[23\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05507__A1 _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10862_ _01291_ io_in[4] u_cpu.rf_ram.memory\[27\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10793_ _01222_ io_in[4] u_cpu.rf_ram.memory\[59\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07680__A1 u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09421__A2 _04605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07983__A2 _03626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05994__A1 _01393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10227_ _00017_ io_in[4] u_cpu.rf_ram_if.rdata1\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08393__C1 _03963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10158_ _00604_ io_in[4] u_cpu.rf_ram.memory\[131\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05746__A1 _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10089_ _00535_ io_in[4] u_cpu.rf_ram.memory\[39\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09488__A2 _04197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[10\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07499__A1 _03353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08696__B1 _04175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09996__D _00003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06320_ _02497_ _02673_ _02677_ _00125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06251_ _02517_ _02628_ _02636_ _00097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06474__A2 _02448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07671__A1 _02311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05202_ _01679_ _01693_ _01694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06182_ _02593_ u_cpu.rf_ram.memory\[1\]\[5\] _02578_ _02594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09412__A2 _04595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10532__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05133_ u_cpu.rf_ram.memory\[32\]\[0\] u_cpu.rf_ram.memory\[33\]\[0\] u_cpu.rf_ram.memory\[34\]\[0\]
+ u_cpu.rf_ram.memory\[35\]\[0\] _01623_ _01624_ _01625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_116_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06226__A2 _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07423__A1 _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07974__A2 _03626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09941_ _00395_ io_in[4] u_cpu.rf_ram.memory\[56\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05064_ _01555_ _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05985__A1 _02305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09176__A1 _04280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09872_ _00326_ io_in[4] u_cpu.rf_ram.memory\[29\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10682__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07726__A2 _03475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08923__A1 _01428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08823_ _03973_ _04256_ _04257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05737__A1 _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08754_ _04211_ _01026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05966_ u_cpu.cpu.state.o_cnt_r\[0\] u_cpu.cpu.state.o_cnt_r\[1\] u_cpu.cpu.state.o_cnt_r\[2\]
+ u_cpu.cpu.state.o_cnt_r\[3\] _02433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_07705_ _03355_ _03465_ _03471_ _00716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04917_ _01437_ u_cpu.cpu.ctrl.o_ibus_adr\[2\] _01439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08685_ _04171_ _00997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_05897_ _02338_ _02378_ _02379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_38_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08151__A2 u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07636_ _03431_ _03432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[28\]_D u_arbiter.i_wb_cpu_rdt\[25\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_04848_ u_cpu.cpu.branch_op _01374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06448__I _02516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05596__S0 _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07567_ u_cpu.rf_ram.memory\[125\]\[1\] _03392_ _03394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08439__B1 _03779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10062__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09306_ _02727_ _04197_ _04535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09100__A1 _04296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06518_ u_cpu.rf_ram.memory\[17\]\[0\] _02801_ _02802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07498_ u_cpu.rf_ram.memory\[22\]\[4\] _03345_ _03354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09237_ _04497_ _01223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07662__A1 _03351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06449_ u_cpu.rf_ram.memory\[50\]\[7\] _02740_ _02755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09168_ _04292_ _04449_ _04455_ _01196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09403__A2 _04595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06217__A2 _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08119_ _03725_ _03678_ _03683_ _03727_ _03728_ _00874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_107_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09099_ u_cpu.rf_ram.memory\[105\]\[7\] _04409_ _04417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07965__A2 _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05976__A1 _01375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08331__C _03876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11061_ _11061_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_1_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08914__A1 _04292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07717__A2 _03475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[33\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10012_ _00458_ io_in[4] u_cpu.rf_ram.memory\[141\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05728__A1 _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05690__C _01628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08678__B1 _04157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10405__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10914_ _01343_ io_in[4] u_cpu.rf_ram.memory\[100\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_u_scanchain_local.scan_flop\[19\]_D u_arbiter.i_wb_cpu_rdt\[16\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08774__S _04217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05587__S0 _01619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10845_ _01274_ io_in[4] u_cpu.rf_ram.memory\[88\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09578__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05900__A1 _01374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05339__S0 _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10776_ _01205_ io_in[4] u_cpu.rf_ram.memory\[69\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10555__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07653__A1 _02561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[61\] u_scanchain_local.module_data_in\[60\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[23\] u_scanchain_local.clk u_scanchain_local.module_data_in\[61\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_12_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05211__B _01565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07405__A1 _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07956__A2 _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05967__A1 _01372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09158__A1 _04280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08949__S _04331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07708__A2 _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05719__A1 _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05820_ u_cpu.cpu.state.o_cnt_r\[0\] u_cpu.cpu.state.o_cnt_r\[1\] u_cpu.cpu.state.o_cnt_r\[2\]
+ u_cpu.cpu.state.o_cnt_r\[3\] _02304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_95_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05751_ _01589_ _02235_ _02236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10085__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08133__A2 _03731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08470_ _03999_ _04028_ _04033_ _04034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05682_ u_cpu.rf_ram.memory\[108\]\[6\] u_cpu.rf_ram.memory\[109\]\[6\] u_cpu.rf_ram.memory\[110\]\[6\]
+ u_cpu.rf_ram.memory\[111\]\[6\] _01598_ _01573_ _02168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_51_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06144__A1 _02492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05578__S0 _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07421_ _03165_ _03305_ _03309_ _00594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07352_ u_cpu.rf_ram.memory\[136\]\[5\] _03265_ _03271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06303_ _02502_ _02662_ _02667_ _00118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07644__A1 _03351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06447__A2 _02740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07283_ _03171_ _03225_ _03232_ _00533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09022_ _04290_ _04369_ _04374_ _01131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06234_ _02625_ _02626_ _02627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05750__S0 _01590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09397__A1 u_cpu.cpu.genblk3.csr.o_new_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06165_ _02580_ _02581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07827__I _02491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07947__A2 _03606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[56\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05116_ _01593_ _01596_ _01600_ _01606_ _01607_ _01608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_46_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06096_ u_cpu.rf_ram.memory\[21\]\[7\] _02530_ _02538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05047_ _01419_ _01420_ _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09924_ _00378_ io_in[4] u_cpu.rf_ram.memory\[58\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09855_ _00309_ io_in[4] u_cpu.rf_ram.memory\[65\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08372__A2 _02313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08806_ _04040_ _04240_ _03780_ _04241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10428__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06383__A1 _02507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06998_ u_cpu.rf_ram.memory\[54\]\[1\] _03071_ _03073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09786_ _00240_ io_in[4] u_cpu.rf_ram.memory\[77\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05186__A2 _01666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08737_ _03545_ _04199_ _04202_ _01018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05949_ _02320_ _02422_ _02423_ _00020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09720__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08124__A2 _03731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09321__A1 _04482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08668_ u_cpu.cpu.ctrl.o_ibus_adr\[5\] _04155_ _04157_ u_cpu.cpu.ctrl.o_ibus_adr\[6\]
+ _04163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06135__A1 _01668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05082__I _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05569__S0 _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10578__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07619_ u_cpu.rf_ram.memory\[38\]\[0\] _03422_ _03423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08599_ u_arbiter.i_wb_cpu_dbus_adr\[20\] u_arbiter.i_wb_cpu_dbus_adr\[19\] _04115_
+ _04122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10630_ _01059_ io_in[4] u_cpu.rf_ram.memory\[97\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09870__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07635__A1 _02524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10561_ _00991_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06438__A2 _02740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10492_ _00925_ io_in[4] u_cpu.cpu.immdec.imm31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05741__S0 _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09388__A1 _02348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07938__A2 _03606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05949__A1 _02320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11113_ u_scanchain_local.clk_out io_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11044_ _11044_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_39_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09560__A1 _03797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08363__A2 _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08115__A2 _02781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06126__A1 _02497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07874__A1 _03549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06677__A2 _02884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10828_ _01257_ io_in[4] u_cpu.rf_ram.memory\[111\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07626__A1 _03351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06429__A2 _02740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10759_ _01188_ io_in[4] u_cpu.rf_ram.memory\[83\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05732__S0 _01546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07929__A2 _03596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08051__A1 u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07970_ _03625_ _03626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06601__A2 _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06921_ _03029_ _00374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09743__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09551__A1 _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08354__A2 _03923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09640_ _00094_ io_in[4] u_cpu.rf_ram.memory\[78\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06852_ _02991_ _02992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_95_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06199__S _02603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05803_ _01609_ _02287_ _02288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09571_ _02783_ _04689_ _01365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06783_ u_cpu.rf_ram.memory\[64\]\[5\] _02944_ _02950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10720__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09303__A1 _04482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08106__A2 _02781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08522_ u_cpu.cpu.genblk3.csr.timer_irq_r _04080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05734_ u_cpu.rf_ram.memory\[12\]\[7\] u_cpu.rf_ram.memory\[13\]\[7\] u_cpu.rf_ram.memory\[14\]\[7\]
+ u_cpu.rf_ram.memory\[15\]\[7\] _01571_ _01668_ _02219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_70_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06117__A1 _02469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09893__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08453_ _04018_ _04016_ _04019_ _03834_ _00917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_63_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05665_ _01540_ _02150_ _01564_ _02151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06668__A2 _02884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06912__I0 _02587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07404_ u_cpu.rf_ram.memory\[133\]\[4\] _03295_ _03300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08384_ _03913_ _03957_ _00910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10870__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05340__A2 _01829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05596_ u_cpu.rf_ram.memory\[104\]\[5\] u_cpu.rf_ram.memory\[105\]\[5\] u_cpu.rf_ram.memory\[106\]\[5\]
+ u_cpu.rf_ram.memory\[107\]\[5\] _01615_ _01616_ _02083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_50_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07617__A1 _02639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07335_ _03169_ _03255_ _03261_ _00556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_17_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07266_ _02599_ u_cpu.rf_ram.memory\[14\]\[7\] _03215_ _03223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07093__A2 _03119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05723__S0 _01680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10100__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09005_ u_cpu.rf_ram.memory\[102\]\[5\] _04359_ _04365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06217_ _02487_ _02614_ _02616_ _00083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05786__B _01626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06840__A2 _02982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07197_ _02602_ _02626_ _03185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04851__A1 u_cpu.cpu.decode.op21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06148_ _02502_ _02563_ _02568_ _00062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06079_ _02527_ _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10250__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08589__S _04115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09907_ _00361_ io_in[4] u_cpu.rf_ram.memory\[19\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08345__A2 _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09542__A1 _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09838_ _00292_ io_in[4] u_cpu.rf_ram.memory\[67\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05159__A2 _01650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06356__A1 _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09769_ _00223_ io_in[4] u_cpu.rf_ram.memory\[129\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06108__A1 _02497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07856__A1 _03549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06659__A2 _02874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05331__A2 _01820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07608__A1 _03351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10613_ _01042_ io_in[4] u_cpu.rf_ram.memory\[93\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09616__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10544_ _00976_ io_in[4] u_cpu.rf_ram.memory\[30\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08281__A1 _03825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07084__A2 _03119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05714__S0 _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05095__A1 _01542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10475_ _00908_ io_in[4] u_cpu.cpu.immdec.imm24_20\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06831__A2 _02972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05190__S1 _01681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04842__A1 u_cpu.cpu.bufreg.lsb\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08033__A1 _02774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09766__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[24\] u_arbiter.i_wb_cpu_rdt\[21\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[18\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_116_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10743__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11027_ _11027_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__09533__A1 _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06347__A1 _02512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06898__A2 _03012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10893__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07147__I0 _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08247__B _03840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05450_ u_cpu.rf_ram.memory\[72\]\[3\] u_cpu.rf_ram.memory\[73\]\[3\] u_cpu.rf_ram.memory\[74\]\[3\]
+ u_cpu.rf_ram.memory\[75\]\[3\] _01610_ _01668_ _01939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05322__A2 _01811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10123__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05381_ _01542_ _01869_ _01870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07120_ u_cpu.rf_ram.memory\[140\]\[0\] _03139_ _03140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08272__A1 _03773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08272__B2 _03755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05705__S0 _01590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07051_ _02581_ u_cpu.rf_ram.memory\[9\]\[1\] _03100_ _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06822__A2 _02972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10273__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05181__S1 _01668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06002_ _02456_ _02458_ _02459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06586__A1 _02750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07953_ u_cpu.rf_ram.memory\[115\]\[0\] _03616_ _03617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09524__A1 _02475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08327__A2 _03860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06904_ _02969_ _03012_ _03020_ _00366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07884_ _02581_ u_cpu.rf_ram.memory\[8\]\[1\] _03577_ _03579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_46_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09623_ _00077_ io_in[4] u_cpu.rf_ram.memory\[7\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06835_ u_cpu.rf_ram.memory\[62\]\[0\] _02982_ _02983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06889__A2 _03012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09554_ u_cpu.rf_ram.memory\[23\]\[5\] _04674_ _04680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06766_ _02750_ _02934_ _02940_ _00308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05561__A2 _02047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05717_ _01553_ _02202_ _01648_ _02203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08505_ u_cpu.cpu.immdec.imm19_12_20\[7\] _04016_ _04066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07838__A1 _03551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09485_ _04641_ _01327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06697_ _02599_ u_cpu.rf_ram.memory\[6\]\[7\] _02894_ _02902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09639__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08436_ _03744_ _03818_ _04004_ _03778_ _04005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05648_ u_cpu.rf_ram.memory\[4\]\[6\] u_cpu.rf_ram.memory\[5\]\[6\] u_cpu.rf_ram.memory\[6\]\[6\]
+ u_cpu.rf_ram.memory\[7\]\[6\] _01578_ _01550_ _02134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__05313__A2 _01802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08367_ _03810_ _03941_ _03763_ _03942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05579_ _01636_ _02065_ _02066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10616__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07318_ u_cpu.rf_ram.memory\[137\]\[6\] _03245_ _03252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08263__A1 _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08298_ _03547_ _03879_ _03883_ _00898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09789__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07249_ u_cpu.rf_ram.memory\[143\]\[7\] _03206_ _03214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06813__A2 _02955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05172__S1 _01652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10260_ _00693_ io_in[4] u_cpu.rf_ram.memory\[37\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08015__A1 u_arbiter.i_wb_cpu_rdt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08015__B2 u_arbiter.i_wb_cpu_dbus_dat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10766__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10191_ _00637_ io_in[4] u_cpu.rf_ram.memory\[128\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09515__A1 _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05552__A2 _02039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10146__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07829__A1 _03545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05304__A2 _01793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06501__A1 _02738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05855__A3 u_cpu.cpu.mem_bytecnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10296__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10527_ _00960_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06804__A2 _02955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08006__A1 u_cpu.cpu.bufreg.lsb\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10458_ _00891_ io_in[4] u_cpu.cpu.csr_d_sel vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08557__A2 _04094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10389_ _00822_ io_in[4] u_cpu.rf_ram.memory\[115\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09506__A1 _02561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05240__A1 _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04950_ u_arbiter.i_wb_cpu_dbus_adr\[8\] _01457_ _01466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08957__S _04331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04881_ u_cpu.cpu.immdec.imm19_12_20\[5\] u_cpu.rf_ram_if.rtrig0 _01407_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_92_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06620_ _02748_ _02854_ _02859_ _00243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05543__A2 _02021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06740__A1 _02742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06551_ u_cpu.rf_ram.memory\[40\]\[7\] _02812_ _02820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05502_ _01541_ _01989_ _01626_ _01990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_33_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09270_ _02625_ _04197_ _04515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10639__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07296__A2 _03235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06482_ _02774_ _02777_ _02778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08493__A1 _03973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08221_ _03769_ _03802_ _03818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05433_ u_cpu.rf_ram.memory\[116\]\[3\] u_cpu.rf_ram.memory\[117\]\[3\] u_cpu.rf_ram.memory\[118\]\[3\]
+ u_cpu.rf_ram.memory\[119\]\[3\] _01623_ _01624_ _01922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_20_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09931__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08152_ _03749_ _03751_ _03752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08245__A1 _03773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07048__A2 _02695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05364_ u_cpu.rf_ram.memory\[76\]\[2\] u_cpu.rf_ram.memory\[77\]\[2\] u_cpu.rf_ram.memory\[78\]\[2\]
+ u_cpu.rf_ram.memory\[79\]\[2\] _01577_ _01549_ _01854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_140_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07103_ _02953_ _03129_ _03130_ _00455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10789__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08796__A2 _04227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08083_ u_arbiter.i_wb_cpu_rdt\[18\] _03669_ _03678_ u_arbiter.i_wb_cpu_dbus_dat\[18\]
+ _03705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05295_ _01554_ _01784_ _01417_ _01785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07034_ u_cpu.rf_ram.memory\[52\]\[1\] _03091_ _03093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08548__A2 _04094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10019__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06559__A1 _02742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07220__A2 _03196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08985_ u_cpu.rf_ram.memory\[101\]\[4\] _04349_ _04354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07936_ _03539_ _03606_ _03607_ _00812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05782__A2 _02266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10169__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07867_ u_cpu.rf_ram.memory\[121\]\[1\] _03568_ _03570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08720__A2 _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09606_ _00060_ io_in[4] u_cpu.rf_ram.memory\[20\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06818_ _02953_ _02972_ _02973_ _00327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_73_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07798_ _03357_ _03520_ _03527_ _00754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09537_ _04480_ _04664_ _04670_ _01350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06749_ u_cpu.rf_ram.memory\[66\]\[6\] _02924_ _02931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05304__B _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08484__A1 _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09468_ _04482_ _04625_ _04632_ _01319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05090__I _01565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08419_ _03788_ _03786_ _03988_ _03899_ _03989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_12_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09399_ _02528_ _02706_ _04594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05393__S1 _01574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07039__A2 _03091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08787__A2 _04227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06798__A1 u_cpu.rf_ram.memory\[29\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05145__S1 _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10312_ _00745_ io_in[4] u_cpu.rf_ram.memory\[35\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08539__A2 _04084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10243_ _00012_ io_in[4] u_cpu.rf_ram_if.rdata0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07211__A2 _03186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10174_ _00620_ io_in[4] u_cpu.rf_ram.memory\[12\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09804__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06722__A1 _02742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09954__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08475__A1 _03779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07278__A2 _03225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10931__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05384__S1 _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05080_ _01571_ _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07450__A2 _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08260__B _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07202__A2 _03186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10311__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08770_ _02584_ u_cpu.rf_ram.memory\[2\]\[2\] _04217_ _04220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05982_ u_arbiter.i_wb_cpu_ibus_adr\[0\] u_cpu.cpu.ctrl.pc_plus_offset_cy_r _02401_
+ _02446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_84_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05175__I _01540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06961__A1 _02953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07721_ _03353_ _03475_ _03480_ _00723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_04933_ u_cpu.cpu.ctrl.o_ibus_adr\[5\] _01451_ _01452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA_u_scanchain_local.scan_flop\[7\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08702__A2 _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07652_ _03359_ _03432_ _03440_ _00694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_04864_ u_cpu.cpu.csr_imm _01390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10461__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05516__A2 _02003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06603_ u_cpu.rf_ram.memory\[139\]\[5\] _02844_ _02850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07583_ u_cpu.rf_ram.memory\[124\]\[0\] _03402_ _03403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09322_ u_cpu.rf_ram.memory\[111\]\[7\] _04536_ _04544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06534_ _02560_ _02637_ _02810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08466__A1 _03835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09253_ _04505_ _04506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06465_ _02763_ _00184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05375__S1 _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08204_ _03767_ _03802_ _03803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05416_ _01422_ _01895_ _01904_ _01905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_09184_ _04290_ _04459_ _04464_ _01203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05778__C _01628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06396_ u_cpu.rf_ram.memory\[48\]\[3\] _02718_ _02722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08135_ _03551_ _03731_ _03737_ _00881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05347_ _01830_ _01832_ _01834_ _01836_ _01607_ _01837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_119_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08066_ u_arbiter.i_wb_cpu_dbus_dat\[13\] _03683_ _03694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07441__A2 _03315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05278_ _01762_ _01764_ _01766_ _01768_ _01568_ _01769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_108_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07017_ _02957_ _03081_ _03083_ _00416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09827__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09194__A2 _04470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[50\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08941__A2 _04322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08968_ _04344_ _01107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08597__S _04115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10804__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05085__I _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05755__A2 _02239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07919_ u_cpu.rf_ram.memory\[112\]\[1\] _03596_ _03598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08899_ u_cpu.rf_ram.memory\[95\]\[7\] _04299_ _04307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09977__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10930_ _01358_ io_in[4] u_cpu.rf_ram.memory\[23\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05507__A2 _01994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06704__A1 _02742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[65\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10861_ _01290_ io_in[4] u_cpu.rf_ram.memory\[27\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10954__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10792_ _01221_ io_in[4] u_cpu.rf_ram.memory\[59\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05969__B _01445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08209__A1 _03765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07432__A2 _03315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10334__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09185__A2 _04459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10226_ _00016_ io_in[4] u_cpu.rf_ram_if.rdata1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07196__A1 _03173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[18\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08393__C2 _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08932__A2 _04322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10157_ _00603_ io_in[4] u_cpu.rf_ram.memory\[131\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10484__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06943__A1 _02953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05746__A2 _02230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10088_ _00534_ io_in[4] u_cpu.rf_ram.memory\[138\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07499__A2 _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08999__A2 _04359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06250_ u_cpu.rf_ram.memory\[78\]\[7\] _02628_ _02636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09248__I0 _02596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07671__A2 _02773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05201_ _01683_ _01686_ _01690_ _01692_ _01404_ _01693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_06181_ _02592_ _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05132_ _01547_ _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07423__A2 _03305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05434__A1 _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05063_ _01543_ _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09940_ _00394_ io_in[4] u_cpu.rf_ram.memory\[56\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10827__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05985__A2 _02448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09176__A2 _04459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09871_ _00325_ io_in[4] u_cpu.rf_ram.memory\[29\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08822_ _03782_ _04255_ _04256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05737__A2 _02221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08753_ _02584_ u_cpu.rf_ram.memory\[3\]\[2\] _04208_ _04211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05965_ _02332_ _02431_ _01409_ _02361_ _02432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_66_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04958__B _01442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07704_ u_cpu.rf_ram.memory\[91\]\[5\] _03465_ _03471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04916_ _01437_ u_cpu.cpu.ctrl.o_ibus_adr\[2\] _01438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_94_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08684_ u_cpu.cpu.ctrl.o_ibus_adr\[13\] _04155_ _04157_ u_cpu.cpu.ctrl.o_ibus_adr\[14\]
+ _04171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05896_ _02376_ u_cpu.cpu.ctrl.i_iscomp _02377_ _02378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_54_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07635_ _02524_ _02639_ _03431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04847_ _01372_ _01373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_26_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10207__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05596__S1 _01616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08439__A1 _03763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07566_ _03343_ _03392_ _03393_ _00655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08439__B2 _03744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09100__A2 _04409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09305_ _04484_ _04526_ _04534_ _01254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06517_ _02800_ _02801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07111__A1 _02963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07497_ _02501_ _03353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09236_ _02573_ u_cpu.rf_ram.memory\[10\]\[0\] _04496_ _04497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07662__A2 _03442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06448_ _02516_ _02754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10357__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09167_ u_cpu.rf_ram.memory\[108\]\[5\] _04449_ _04455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06379_ _02497_ _02708_ _02712_ _00149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08118_ u_arbiter.i_wb_cpu_rdt\[30\] _02781_ _03728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08072__C1 _03676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07414__A2 _03305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09098_ _04294_ _04409_ _04416_ _01165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05425__A1 _01601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08049_ _03682_ _00850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_135_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05976__A2 _02356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11060_ _11060_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__09167__A2 _04449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07178__A1 _03173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10011_ _00457_ io_in[4] u_cpu.rf_ram.memory\[141\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08914__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05728__A2 _02213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06925__A1 _02953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10913_ _01342_ io_in[4] u_cpu.rf_ram.memory\[100\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06153__A2 _02563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05587__S1 _01620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10844_ _01273_ io_in[4] u_cpu.rf_ram.memory\[88\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09478__I0 _02587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05900__A2 _02313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10775_ _01204_ io_in[4] u_cpu.rf_ram.memory\[69\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05339__S1 _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08850__A1 _03549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07653__A2 _02639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[54\] u_scanchain_local.module_data_in\[53\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[16\] u_scanchain_local.clk u_scanchain_local.module_data_in\[54\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_126_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07405__A2 _03295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05416__A1 _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06464__I0 _02596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05967__A2 _01374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09158__A2 _04449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07169__A1 _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08905__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10209_ _00655_ io_in[4] u_cpu.rf_ram.memory\[125\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05719__A2 _02195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06392__A2 _02718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05750_ u_cpu.rf_ram.memory\[52\]\[7\] u_cpu.rf_ram.memory\[53\]\[7\] u_cpu.rf_ram.memory\[54\]\[7\]
+ u_cpu.rf_ram.memory\[55\]\[7\] _01590_ _01591_ _02235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08965__S _04331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09330__A2 _04546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05681_ _01539_ _02138_ _02147_ _02166_ _02167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_36_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06144__A2 _02563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05578__S1 _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07420_ u_cpu.rf_ram.memory\[132\]\[3\] _03305_ _03309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07351_ _03167_ _03265_ _03270_ _00563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09094__A1 _04290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08141__I0 u_arbiter.i_wb_cpu_rdt\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06302_ u_cpu.rf_ram.memory\[45\]\[4\] _02662_ _02667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09672__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07282_ u_cpu.rf_ram.memory\[138\]\[6\] _03225_ _03232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07644__A2 _03432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09021_ u_cpu.rf_ram.memory\[103\]\[4\] _04369_ _04374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06233_ _02473_ _02575_ _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05750__S1 _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06164_ u_cpu.rf_ram_if.wdata0_r\[1\] u_cpu.rf_ram_if.wdata1_r\[1\] _02478_ _02580_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09397__A2 _03458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05115_ _01425_ _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06095_ _02512_ _02530_ _02537_ _00040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05958__A2 _01403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06080__A1 _02524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09149__A2 _04439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05046_ _01538_ u_arbiter.o_wb_cpu_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09923_ _00377_ io_in[4] u_cpu.rf_ram.memory\[58\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06207__I0 _02596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09854_ _00308_ io_in[4] u_cpu.rf_ram.memory\[65\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08805_ _03857_ _03897_ _04239_ _04240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09785_ _00239_ io_in[4] u_cpu.rf_ram.memory\[77\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07580__A1 _03359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06383__A2 _02708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08109__B1 _03654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06997_ _02953_ _03071_ _03072_ _00407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05186__A3 _01677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08736_ u_cpu.rf_ram.memory\[109\]\[2\] _04199_ _04202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05948_ _02320_ u_cpu.rf_ram_if.rdata1\[6\] _02423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09321__A2 _04536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08667_ _04162_ _00988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05879_ u_cpu.cpu.bufreg.lsb\[0\] _02361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_54_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05569__S1 _01574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07618_ _03421_ _03422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_81_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08598_ _04121_ _00960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07549_ u_cpu.rf_ram.memory\[126\]\[1\] _03382_ _03384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07635__A2 _02639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10560_ _00990_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09219_ u_cpu.rf_ram.memory\[59\]\[0\] _04487_ _04488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10491_ _00924_ io_in[4] u_cpu.cpu.immdec.imm19_12_20\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05741__S1 _01574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07399__A1 _03161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08060__A2 _03683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06071__A1 _01547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11112_ io_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_1_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11043_ _11043_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_122_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05257__S0 _01623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09560__A2 _03458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06374__A2 _02708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09312__A2 _04536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10522__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06126__A2 _02551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08520__B1 _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09695__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07874__A2 _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05885__A1 _01373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10827_ _01256_ io_in[4] u_cpu.rf_ram.memory\[111\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09076__A1 _04290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10672__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10758_ _01187_ io_in[4] u_cpu.rf_ram.memory\[83\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07626__A2 _03422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08823__A1 _03973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06685__I0 _02581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10689_ _01118_ io_in[4] u_cpu.rf_ram.memory\[101\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05732__S1 _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08051__A2 _03683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06920_ _02599_ u_cpu.rf_ram.memory\[5\]\[7\] _03021_ _03029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10052__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09000__A1 _04286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05248__S0 _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09551__A2 _04674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06851_ _02660_ _02684_ _02991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07562__A1 _03359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06365__A2 _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05802_ u_cpu.rf_ram.memory\[72\]\[7\] u_cpu.rf_ram.memory\[73\]\[7\] u_cpu.rf_ram.memory\[74\]\[7\]
+ u_cpu.rf_ram.memory\[75\]\[7\] _01610_ _01611_ _02287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09570_ _02769_ _04688_ _04689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06782_ _02748_ _02944_ _02949_ _00315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09303__A2 _04526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08521_ _03798_ _03906_ _04077_ _04079_ _00925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_82_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05733_ _01542_ _02217_ _02218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05116__C _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06117__A2 _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08452_ u_cpu.cpu.immdec.imm19_12_20\[2\] _03797_ _04016_ _04019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_35_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07865__A2 _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05664_ u_cpu.rf_ram.memory\[48\]\[6\] u_cpu.rf_ram.memory\[49\]\[6\] u_cpu.rf_ram.memory\[50\]\[6\]
+ u_cpu.rf_ram.memory\[51\]\[6\] _01544_ _01548_ _02150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__05420__S0 _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05876__A1 _02309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07403_ _03165_ _03295_ _03299_ _00586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_91_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05595_ _01597_ _02081_ _02082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08383_ u_cpu.cpu.immdec.imm30_25\[1\] _03954_ _03956_ u_cpu.cpu.immdec.imm30_25\[2\]
+ _03957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_91_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07334_ u_cpu.rf_ram.memory\[49\]\[5\] _03255_ _03261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07617__A2 _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[23\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08814__A1 _03762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07265_ _03222_ _00525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09004_ _04290_ _04359_ _04364_ _01123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05723__S1 _01681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06216_ u_cpu.rf_ram.memory\[80\]\[1\] _02614_ _02616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07196_ _03173_ _03176_ _03184_ _00494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06147_ u_cpu.rf_ram.memory\[20\]\[4\] _02563_ _02568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06053__A1 _02460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06078_ u_cpu.cpu.immdec.imm11_7\[3\] _02470_ _02526_ _02527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_132_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05029_ _01445_ _01524_ _01525_ u_arbiter.o_wb_cpu_adr\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_59_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09906_ _00360_ io_in[4] u_cpu.rf_ram.memory\[19\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09542__A2 _02602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09837_ _00291_ io_in[4] u_cpu.rf_ram.memory\[67\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10545__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06356__A2 _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[30\]_SI u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09768_ _00222_ io_in[4] u_cpu.rf_ram.memory\[119\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08719_ _04189_ _01013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_73_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06108__A2 _02541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09699_ _00153_ io_in[4] u_cpu.rf_ram.memory\[43\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10695__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07856__A2 _03558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05867__A1 u_arbiter.i_wb_cpu_ibus_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05411__S0 _01619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09058__A1 _04290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10612_ _01041_ io_in[4] u_cpu.rf_ram.memory\[93\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07608__A2 _03412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10543_ _00975_ io_in[4] u_cpu.cpu.bufreg.lsb\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05714__S1 _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06292__A1 _02639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05095__A2 _01586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10474_ _00907_ io_in[4] u_cpu.cpu.immdec.imm24_20\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04842__A2 u_cpu.cpu.bufreg.lsb\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10075__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09230__A1 _04480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07792__A1 _03351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06595__A2 _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[17\] u_arbiter.i_wb_cpu_rdt\[14\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[11\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_89_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07483__I _02481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11026_ _11026_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__09533__A2 _04664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04900__I _01425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07544__A1 _03359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06347__A2 _02686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05650__S0 _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09297__A1 _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07847__A2 _03558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[46\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05402__S0 _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05380_ u_cpu.rf_ram.memory\[8\]\[3\] u_cpu.rf_ram.memory\[9\]\[3\] u_cpu.rf_ram.memory\[10\]\[3\]
+ u_cpu.rf_ram.memory\[11\]\[3\] _01546_ _01550_ _01869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_118_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08272__A2 _03860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05705__S1 _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10418__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08263__B _03854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07050_ _03101_ _00431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_12_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06001_ _02312_ _02457_ _02458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09710__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08024__A2 _02774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06035__A1 _02460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10568__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07783__A1 _02469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06586__A2 _02834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07952_ _03615_ _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09524__A2 _02695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06903_ u_cpu.rf_ram.memory\[19\]\[7\] _03012_ _03020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09860__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07883_ _03578_ _00788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06338__A2 _02686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09622_ _00076_ io_in[4] u_cpu.rf_ram.memory\[7\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06834_ _02981_ _02982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09553_ _04478_ _04674_ _04679_ _01357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09288__A1 _02475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06765_ u_cpu.rf_ram.memory\[65\]\[5\] _02934_ _02940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08504_ u_cpu.cpu.immdec.imm19_12_20\[8\] _02768_ _04065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_70_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05716_ u_cpu.rf_ram.memory\[76\]\[6\] u_cpu.rf_ram.memory\[77\]\[6\] u_cpu.rf_ram.memory\[78\]\[6\]
+ u_cpu.rf_ram.memory\[79\]\[6\] _01577_ _01549_ _02202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_93_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07838__A2 _03541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09484_ _02596_ u_cpu.rf_ram.memory\[0\]\[6\] _04634_ _04641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06696_ _02901_ _00277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08435_ _03999_ _03776_ _04004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05647_ _01554_ _02132_ _01417_ _02133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06510__A2 _02791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08366_ _03785_ _03891_ _03941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05578_ u_cpu.rf_ram.memory\[60\]\[5\] u_cpu.rf_ram.memory\[61\]\[5\] u_cpu.rf_ram.memory\[62\]\[5\]
+ u_cpu.rf_ram.memory\[63\]\[5\] _01598_ _01573_ _02065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_108_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07317_ _03169_ _03245_ _03251_ _00548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10098__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08297_ u_cpu.rf_ram.memory\[114\]\[3\] _03879_ _03883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09460__A1 _04474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07248_ _03171_ _03206_ _03213_ _00517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08015__A2 _03653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07179_ _02626_ _02695_ _03175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05088__I _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07074__I0 _02590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10190_ _00636_ io_in[4] u_cpu.rf_ram.memory\[128\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07774__A1 _03351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06577__A2 _02834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09515__A2 _04654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07526__A1 _03359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[69\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09279__A1 _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08348__B _03759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07829__A2 _03541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06501__A2 _02791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08862__I _02486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09733__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10526_ _00959_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10710__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08006__A2 u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10457_ _00890_ io_in[4] u_cpu.cpu.decode.co_mem_word vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06017__A1 u_cpu.cpu.immdec.imm11_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09883__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10388_ _00821_ io_in[4] u_cpu.rf_ram.memory\[115\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07765__A1 _02639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06568__A2 _02823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10860__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09506__A2 _04197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08714__B1 _04175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11009_ _11009_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_04880_ _01405_ _01406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08190__A1 _03785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05543__A3 _02030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06740__A2 _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06550_ _02752_ _02812_ _02819_ _00213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_46_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08973__S _04331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05501_ u_cpu.rf_ram.memory\[32\]\[4\] u_cpu.rf_ram.memory\[33\]\[4\] u_cpu.rf_ram.memory\[34\]\[4\]
+ u_cpu.rf_ram.memory\[35\]\[4\] _01623_ _01624_ _01989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_34_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06481_ u_arbiter.i_wb_cpu_dbus_dat\[5\] _02776_ _02777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08220_ _03814_ _03817_ _00886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10240__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05432_ _01541_ _01920_ _01921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08151_ _02765_ u_arbiter.i_wb_cpu_rdt\[12\] _03750_ _03751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10954__D u_cpu.cpu.o_wdata1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05363_ _01667_ _01852_ _01853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08245__A2 _03767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09442__A1 _04474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07102_ u_cpu.rf_ram.memory\[141\]\[0\] _03129_ _03130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05410__B _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05294_ u_cpu.rf_ram.memory\[12\]\[2\] u_cpu.rf_ram.memory\[13\]\[2\] u_cpu.rf_ram.memory\[14\]\[2\]
+ u_cpu.rf_ram.memory\[15\]\[2\] _01556_ _01557_ _01784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08082_ u_arbiter.i_wb_cpu_dbus_dat\[19\] _03683_ _03704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10390__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07033_ _02953_ _03091_ _03092_ _00423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07756__A1 _03351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06559__A2 _02823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08984_ _04288_ _04349_ _04353_ _01114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07935_ u_cpu.rf_ram.memory\[122\]\[0\] _03606_ _03607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07508__A1 _03359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07866_ _03539_ _03568_ _03569_ _00780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09606__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08181__A1 _03779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09605_ _00059_ io_in[4] u_cpu.rf_ram.memory\[20\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06817_ u_cpu.rf_ram.memory\[63\]\[0\] _02972_ _02973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07797_ u_cpu.rf_ram.memory\[34\]\[6\] _03520_ _03527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06731__A2 _02914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09536_ u_cpu.rf_ram.memory\[89\]\[5\] _04664_ _04670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06748_ _02750_ _02924_ _02930_ _00300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09756__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09467_ u_cpu.rf_ram.memory\[24\]\[6\] _04625_ _04632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06679_ u_cpu.rf_ram.memory\[75\]\[7\] _02884_ _02892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08418_ _03802_ _03826_ _03988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_40_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09398_ _01428_ u_cpu.cpu.genblk3.csr.timer_irq_r _04082_ _04593_ _01288_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_8_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10733__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08349_ _03871_ _03925_ _03926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06247__A1 _02507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06798__A2 _02955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10311_ _00744_ io_in[4] u_cpu.rf_ram.memory\[35\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10883__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10242_ _00011_ io_in[4] u_cpu.rf_ram_if.rdata0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07747__A1 _02475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10173_ _00619_ io_in[4] u_cpu.rf_ram.memory\[12\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10113__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06970__A2 _03051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08857__I _02481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04981__A1 _01443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05605__S0 _01646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06722__A2 _02914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10263__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08806__B _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06486__A1 _01373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09424__A1 _04474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07986__A1 _03555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10509_ _00942_ io_in[4] u_cpu.rf_ram.memory\[31\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09629__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06410__A1 _02482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05981_ _02439_ _02444_ _02445_ _00022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06961__A2 _03051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07720_ u_cpu.rf_ram.memory\[90\]\[4\] _03475_ _03480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04932_ _01434_ u_cpu.cpu.ctrl.o_ibus_adr\[4\] u_cpu.cpu.ctrl.o_ibus_adr\[3\] u_cpu.cpu.ctrl.o_ibus_adr\[2\]
+ _01451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__10606__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04972__A1 _01443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07651_ u_cpu.rf_ram.memory\[37\]\[7\] _03432_ _03440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04863_ u_cpu.cpu.immdec.imm24_20\[0\] _01388_ _01389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09779__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06713__A2 _02904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06602_ _02748_ _02844_ _02849_ _00235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05405__B _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07582_ _03401_ _03402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_92_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09321_ _04482_ _04536_ _04543_ _01261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10756__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06533_ _02754_ _02801_ _02809_ _00206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08466__A2 _03988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09252_ _02475_ _02524_ _04505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06464_ _02596_ u_cpu.rf_ram.memory\[4\]\[6\] _02756_ _02763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_138_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08203_ u_arbiter.i_wb_cpu_rdt\[13\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[13\]
+ _01436_ _03802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05415_ _01897_ _01899_ _01901_ _01903_ _01628_ _01904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_09183_ u_cpu.rf_ram.memory\[69\]\[4\] _04459_ _04464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06395_ _02492_ _02718_ _02721_ _00156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06229__A1 _02517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08134_ u_cpu.rf_ram.memory\[113\]\[5\] _03731_ _03737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05346_ _01614_ _01835_ _01654_ _01836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_105_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08065_ _03692_ _03693_ _00855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05277_ _01636_ _01767_ _01417_ _01768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_108_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07016_ u_cpu.rf_ram.memory\[53\]\[1\] _03081_ _03083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10136__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07729__A1 u_cpu.cpu.state.genblk1.misalign_trap_sync_r vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06401__A1 _02507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08967_ u_arbiter.i_wb_cpu_rdt\[28\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[12\]
+ _04331_ _04344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_76_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06952__A2 _03041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10286__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07918_ _03539_ _03596_ _03597_ _00804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08898_ _04294_ _04299_ _04306_ _01075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08154__A1 _02765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07849_ u_cpu.rf_ram.memory\[118\]\[1\] _03558_ _03560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06704__A2 _02904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10860_ _01289_ io_in[4] u_cpu.rf_ram.memory\[27\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09519_ _04480_ _04654_ _04660_ _01342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08457__A2 _04016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10791_ _01220_ io_in[4] u_cpu.rf_ram.memory\[59\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08209__A2 _03778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09406__A1 _04474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07968__A1 _03555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06640__A1 _02750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08768__I0 _02581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10225_ _00015_ io_in[4] u_cpu.rf_ram_if.rdata1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10629__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07196__A2 _03176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10156_ _00602_ io_in[4] u_cpu.rf_ram.memory\[131\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06943__A2 _03041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09921__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04954__A1 _01445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10087_ _00533_ io_in[4] u_cpu.rf_ram.memory\[138\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08145__A1 _03741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07491__I _02491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10779__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08696__A2 _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05225__B _01564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05903__B1 u_cpu.cpu.mem_bytecnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10989_ _10989_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_43_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10009__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09211__I _02511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07120__A2 _03139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08255__C _03800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05200_ _01684_ _01691_ _01418_ _01692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06180_ u_cpu.rf_ram_if.wdata0_r\[5\] u_cpu.rf_ram_if.wdata1_r\[5\] _02478_ _02592_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10159__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05131_ _01544_ _01623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05062_ _01553_ _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08759__I0 _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09870_ _00324_ io_in[4] u_cpu.rf_ram.memory\[29\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08384__A1 _03913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07187__A2 _03176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08821_ _03825_ _03770_ _04255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05198__A1 _01399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06934__A2 _03031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08752_ _04210_ _01025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05964_ u_cpu.cpu.bufreg.lsb\[1\] _02431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_39_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07703_ _03353_ _03465_ _03470_ _00715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04915_ _01436_ _01437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_54_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08683_ _04170_ _00996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_66_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05895_ u_cpu.cpu.state.o_cnt_r\[2\] u_cpu.cpu.ctrl.i_iscomp _02377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05135__B _01626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07634_ _03359_ _03422_ _03430_ _00686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_93_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04846_ u_cpu.cpu.decode.opcode\[2\] _01372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07565_ u_cpu.rf_ram.memory\[125\]\[0\] _03392_ _03393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05370__A1 _01399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08439__A2 _03778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__04974__B _01442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09304_ u_cpu.rf_ram.memory\[86\]\[7\] _04526_ _04534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06516_ _02528_ _02539_ _02800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07496_ _03351_ _03345_ _03352_ _00626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07111__A2 _03129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09235_ _02577_ _02638_ _04496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06447_ _02752_ _02740_ _02753_ _00176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06170__I0 _02584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09166_ _04290_ _04449_ _04454_ _01195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06378_ u_cpu.rf_ram.memory\[43\]\[3\] _02708_ _02712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08117_ u_arbiter.i_wb_cpu_dbus_dat\[31\] _03727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08072__B1 _03654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05329_ _01539_ _01790_ _01799_ _01818_ _01819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_09097_ u_cpu.rf_ram.memory\[105\]\[6\] _04409_ _04416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06622__A1 _02750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08048_ u_arbiter.i_wb_cpu_rdt\[6\] _03653_ _03654_ u_arbiter.i_wb_cpu_dbus_dat\[6\]
+ _03676_ u_arbiter.i_wb_cpu_dbus_dat\[7\] _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_134_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09944__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07178__A2 _03159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08375__A1 _02765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10010_ _00456_ io_in[4] u_cpu.rf_ram.memory\[141\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09999_ _00006_ io_in[4] u_cpu.rf_ram.rdata\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10921__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06925__A2 _03031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08127__A1 _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08678__A2 _04155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10912_ _01341_ io_in[4] u_cpu.rf_ram.memory\[100\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07350__A2 _03265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10843_ _01272_ io_in[4] u_cpu.rf_ram.memory\[88\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05361__A1 _01553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05699__C _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10774_ _01203_ io_in[4] u_cpu.rf_ram.memory\[69\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07102__A2 _03129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10301__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08850__A2 _04271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[47\] u_scanchain_local.module_data_in\[46\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[9\] u_scanchain_local.clk u_scanchain_local.module_data_in\[47\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__10451__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__04903__I _01403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07169__A2 _03159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08366__A1 _03785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10208_ _00654_ io_in[4] u_cpu.rf_ram.memory\[126\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05719__A3 _02204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04927__A1 _01445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.input_buf_clk_I io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10139_ _00585_ io_in[4] u_cpu.rf_ram.memory\[133\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08118__A1 u_arbiter.i_wb_cpu_rdt\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05680_ _01422_ _02156_ _02165_ _02166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_39_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05352__A1 _01645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07350_ u_cpu.rf_ram.memory\[136\]\[4\] _03265_ _03270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09817__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09094__A2 _04409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06301_ _02497_ _02662_ _02666_ _00117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07281_ _03169_ _03225_ _03231_ _00532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05104__A1 _01594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08841__A2 _04271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09020_ _04288_ _04369_ _04373_ _01130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06232_ _02468_ _02624_ _02625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_15_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06163_ _02579_ _00066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09967__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06604__A1 _02750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05114_ _01601_ _01604_ _01605_ _01606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_u_scanchain_local.scan_flop\[64\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06094_ u_cpu.rf_ram.memory\[21\]\[6\] _02530_ _02537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10944__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05045_ u_arbiter.i_wb_cpu_dbus_adr\[31\] _01537_ _01431_ _01538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09922_ _00376_ io_in[4] u_cpu.rf_ram.memory\[58\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06080__A2 _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08357__A1 _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09853_ _00307_ io_in[4] u_cpu.rf_ram.memory\[65\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08804_ _03860_ _03818_ _03788_ _04239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04918__A1 _01431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09784_ _00238_ io_in[4] u_cpu.rf_ram.memory\[139\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08109__A1 u_arbiter.i_wb_cpu_rdt\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06996_ u_cpu.rf_ram.memory\[54\]\[0\] _03071_ _03072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07580__A2 _03392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08735_ _03543_ _04199_ _04201_ _01017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05947_ _02321_ u_cpu.rf_ram.rdata\[6\] _02422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05591__B2 _02077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08666_ u_cpu.cpu.ctrl.o_ibus_adr\[4\] _04155_ _04157_ u_cpu.cpu.ctrl.o_ibus_adr\[5\]
+ _04162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05878_ _01410_ _02359_ _02360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07332__A2 _03255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10324__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07617_ _02639_ _02893_ _03421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08597_ u_arbiter.i_wb_cpu_dbus_adr\[19\] u_arbiter.i_wb_cpu_dbus_adr\[18\] _04115_
+ _04121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_54_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07548_ _03343_ _03382_ _03383_ _00647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09085__A2 _04409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[17\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07479_ _02596_ u_cpu.rf_ram.memory\[12\]\[6\] _03334_ _03341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10474__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09218_ _04486_ _04487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10490_ _00923_ io_in[4] u_cpu.cpu.immdec.imm19_12_20\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09149_ u_cpu.rf_ram.memory\[83\]\[5\] _04439_ _04445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07399__A2 _03295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11111_ io_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_2_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11042_ _11042_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_110_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08899__A2 _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05257__S1 _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07571__A2 _03392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08865__I _02491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08520__A1 u_cpu.cpu.immdec.imm31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08520__B2 _04078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10826_ _01255_ io_in[4] u_cpu.rf_ram.memory\[111\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05885__A2 _01370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10817__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09076__A2 _04399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07087__A1 _02957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10757_ _01186_ io_in[4] u_cpu.rf_ram.memory\[83\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08284__B1 _03779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07882__I0 _02573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10688_ _01117_ io_in[4] u_cpu.rf_ram.memory\[101\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05193__S0 _01680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06062__A2 _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08339__A1 _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09000__A2 _04359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07011__A1 _02969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05248__S1 _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06850_ _02969_ _02982_ _02990_ _00342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07562__A2 _03382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05801_ _01553_ _02285_ _01654_ _02286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10347__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06781_ u_cpu.rf_ram.memory\[64\]\[4\] _02944_ _02949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08520_ u_cpu.cpu.immdec.imm31 _03798_ _03816_ _04078_ _04079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_64_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09380__B _01386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05732_ u_cpu.rf_ram.memory\[8\]\[7\] u_cpu.rf_ram.memory\[9\]\[7\] u_cpu.rf_ram.memory\[10\]\[7\]
+ u_cpu.rf_ram.memory\[11\]\[7\] _01546_ _01550_ _02217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_64_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08511__A1 _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07314__A2 _03245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08451_ u_cpu.cpu.immdec.imm19_12_20\[1\] _04018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05663_ _01589_ _02148_ _02149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10497__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07402_ u_cpu.rf_ram.memory\[133\]\[3\] _03295_ _03299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05420__S1 _01616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08382_ _02768_ _03948_ _03956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05594_ u_cpu.rf_ram.memory\[108\]\[5\] u_cpu.rf_ram.memory\[109\]\[5\] u_cpu.rf_ram.memory\[110\]\[5\]
+ u_cpu.rf_ram.memory\[111\]\[5\] _01598_ _01573_ _02081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09067__A2 _04399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07333_ _03167_ _03255_ _03260_ _00555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08814__A2 _03778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07264_ _02596_ u_cpu.rf_ram.memory\[14\]\[6\] _03215_ _03222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09003_ u_cpu.rf_ram.memory\[102\]\[4\] _04359_ _04364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06215_ _02482_ _02614_ _02615_ _00082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07195_ u_cpu.rf_ram.memory\[73\]\[7\] _03176_ _03184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06146_ _02497_ _02563_ _02567_ _00061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07250__A1 _03173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06077_ _02525_ _02472_ _02526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05028_ u_arbiter.i_wb_cpu_dbus_adr\[27\] _01457_ _01525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09905_ _00359_ io_in[4] u_cpu.rf_ram.memory\[19\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09836_ _00290_ io_in[4] u_cpu.rf_ram.memory\[67\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07553__A2 _03382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09767_ _00221_ io_in[4] u_cpu.rf_ram.memory\[119\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06979_ _02953_ _03061_ _03062_ _00399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_73_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08718_ u_cpu.cpu.ctrl.o_ibus_adr\[29\] _04173_ _04175_ u_cpu.cpu.ctrl.o_ibus_adr\[30\]
+ _04189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_73_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09698_ _00152_ io_in[4] u_cpu.rf_ram.memory\[43\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08649_ _03551_ _04145_ _04151_ _00981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05411__S1 _01620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05867__A2 _01386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09058__A2 _04389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10611_ _01040_ io_in[4] u_cpu.rf_ram.memory\[93\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08805__A2 _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10542_ _00974_ io_in[4] u_cpu.cpu.bufreg.lsb\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08353__C _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06292__A2 _02660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10473_ _00906_ io_in[4] u_cpu.cpu.immdec.imm24_20\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09230__A2 _04487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06044__A2 _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05993__B _02453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07792__A2 _03520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11025_ _11025_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_77_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08741__A1 _03549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07544__A2 _03372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09662__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05555__A1 _01406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05650__S1 _01557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09297__A2 _04526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05402__S1 _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09049__A2 _04389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10809_ _01238_ io_in[4] u_cpu.rf_ram.memory\[85\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06807__A1 u_cpu.rf_ram.memory\[29\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05166__S0 _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06283__A2 _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06000_ u_cpu.rf_ram_if.genblk1.wtrig0_r _01386_ _02457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_126_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09221__A2 _04487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07232__A1 _03173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07783__A2 _02639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08980__A1 _04284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07951_ _02682_ _02821_ _03615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05794__A1 _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06902_ _02967_ _03012_ _03019_ _00365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07882_ _02573_ u_cpu.rf_ram.memory\[8\]\[0\] _03577_ _03578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07535__A2 _03372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09621_ _00075_ io_in[4] u_cpu.rf_ram.memory\[7\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06833_ _02625_ _02684_ _02981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05546__A1 _01399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09552_ u_cpu.rf_ram.memory\[23\]\[4\] _04674_ _04679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06764_ _02748_ _02934_ _02939_ _00307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09288__A2 _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08503_ _03782_ _04059_ _04063_ _03797_ _04064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_102_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05715_ _01667_ _02200_ _02201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07299__A1 _03169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09483_ _04640_ _01326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06695_ _02596_ u_cpu.rf_ram.memory\[6\]\[6\] _02894_ _02901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_36_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05143__B _01416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08434_ _03831_ _03828_ _04003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05646_ u_cpu.rf_ram.memory\[12\]\[6\] u_cpu.rf_ram.memory\[13\]\[6\] u_cpu.rf_ram.memory\[14\]\[6\]
+ u_cpu.rf_ram.memory\[15\]\[6\] _01571_ _01557_ _02132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_24_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08365_ _03773_ _03767_ _03940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05577_ _01540_ _02063_ _01564_ _02064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08799__A1 _03555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07316_ u_cpu.rf_ram.memory\[137\]\[5\] _03245_ _03251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08296_ _03545_ _03879_ _03882_ _00897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05797__C _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09460__A2 _04625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07247_ u_cpu.rf_ram.memory\[143\]\[6\] _03206_ _03213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07178_ _03173_ _03159_ _03174_ _00486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_127_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09212__A2 _04470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10512__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06026__A2 _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06129_ u_cpu.rf_ram.memory\[18\]\[5\] _02551_ _02557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07774__A2 _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09685__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10662__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08723__A1 _04191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07526__A2 _03362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09819_ _00273_ io_in[4] u_cpu.rf_ram.memory\[6\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05537__A1 _01553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09279__A2 _04516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09240__S _04496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10042__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09451__A2 _04615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06265__A2 _02641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10525_ _00958_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[7\]_D u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10456_ _00889_ io_in[4] u_cpu.cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09203__A2 _04470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10192__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07214__A1 _03173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10387_ _00820_ io_in[4] u_cpu.rf_ram.memory\[115\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07494__I _02496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07765__A2 _02682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05240__A3 _01730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[13\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07517__A2 _03362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11008_ _11008_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_37_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05528__A1 _01645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09214__I _02516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05500_ _01589_ _01987_ _01988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06480_ u_arbiter.i_wb_cpu_dbus_dat\[4\] _02775_ _02776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05431_ u_cpu.rf_ram.memory\[112\]\[3\] u_cpu.rf_ram.memory\[113\]\[3\] u_cpu.rf_ram.memory\[114\]\[3\]
+ u_cpu.rf_ram.memory\[115\]\[3\] _01619_ _01620_ _01920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_20_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05700__A1 _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08150_ _01436_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[12\] _03750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_119_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05362_ u_cpu.rf_ram.memory\[72\]\[2\] u_cpu.rf_ram.memory\[73\]\[2\] u_cpu.rf_ram.memory\[74\]\[2\]
+ u_cpu.rf_ram.memory\[75\]\[2\] _01571_ _01668_ _01852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA_u_scanchain_local.out_flop_CLKN u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09442__A2 _04615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07101_ _03128_ _03129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10535__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[20\]_SI u_arbiter.i_wb_cpu_dbus_dat\[14\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08081_ _03703_ _00861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__07453__A1 _03161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05293_ _01542_ _01782_ _01783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05189__I _01668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07032_ u_cpu.rf_ram.memory\[52\]\[0\] _03091_ _03092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10685__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07756__A2 _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08983_ u_cpu.rf_ram.memory\[101\]\[3\] _04349_ _04353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05767__B2 _02251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07934_ _03605_ _03606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07508__A2 _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07865_ u_cpu.rf_ram.memory\[121\]\[0\] _03568_ _03569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04977__B u_cpu.cpu.ctrl.o_ibus_adr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08449__B _04016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08181__A2 _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09604_ _00058_ io_in[4] u_cpu.rf_ram.memory\[20\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06816_ _02971_ _02972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07796_ _03355_ _03520_ _03526_ _00753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09535_ _04478_ _04664_ _04669_ _01349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06747_ u_cpu.rf_ram.memory\[66\]\[5\] _02924_ _02930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09130__A1 _04290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10065__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09466_ _04480_ _04625_ _04631_ _01318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06678_ _02752_ _02884_ _02891_ _00269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07692__A1 _02475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08417_ _03741_ _03742_ _03841_ _03986_ _03818_ _03987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_05629_ _01553_ _02115_ _01417_ _02116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_106_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09397_ u_cpu.cpu.genblk3.csr.o_new_irq _03458_ _04593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05601__B _01626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08348_ _03870_ _03924_ _03759_ _03925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09433__A2 _04605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06247__A2 _02628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08279_ _03858_ _03862_ _03869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05099__I _01548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10310_ _00743_ io_in[4] u_cpu.rf_ram.memory\[35\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07995__A2 _03636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10241_ _00010_ io_in[4] u_cpu.rf_ram_if.rdata0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07747__A2 _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[36\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10172_ _00618_ io_in[4] u_cpu.rf_ram.memory\[12\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05758__B2 _02242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04887__B u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05605__S1 _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10408__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05930__A1 _01386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09700__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05369__S0 _01680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10558__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07683__A1 u_cpu.cpu.state.o_cnt_r\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09850__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09424__A2 _04605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07435__A1 _03161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06238__A2 _02628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05230__C _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07986__A2 _03626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10508_ _00941_ io_in[4] u_cpu.rf_ram.memory\[31\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05997__A1 u_cpu.cpu.bufreg.lsb\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09188__A1 _04294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08235__I0 u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10439_ _00872_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07738__A2 _02356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08935__A1 _04290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06410__A2 _02729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05980_ _02372_ _02445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04931_ _01445_ _01449_ _01450_ u_arbiter.o_wb_cpu_adr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09360__A1 _02311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10088__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07650_ _03357_ _03432_ _03439_ _00693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_93_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04862_ u_cpu.rf_ram_if.rtrig0 _01377_ _01387_ _01388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_66_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06601_ u_cpu.rf_ram.memory\[139\]\[4\] _02844_ _02849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07581_ _02671_ _02821_ _03401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05921__A1 u_arbiter.i_wb_cpu_ibus_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09112__A1 _04290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09320_ u_cpu.rf_ram.memory\[111\]\[6\] _04536_ _04543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06532_ u_cpu.rf_ram.memory\[17\]\[7\] _02801_ _02809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09251_ _04504_ _01230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06463_ _02762_ _00183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08202_ _03773_ _03800_ _03801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05414_ _01541_ _01902_ _01626_ _01903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05421__B _01416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09182_ _04288_ _04459_ _04463_ _01202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06394_ u_cpu.rf_ram.memory\[48\]\[2\] _02718_ _02721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09415__A2 _04595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08133_ _03549_ _03731_ _03736_ _00880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05345_ u_cpu.rf_ram.memory\[116\]\[2\] u_cpu.rf_ram.memory\[117\]\[2\] u_cpu.rf_ram.memory\[118\]\[2\]
+ u_cpu.rf_ram.memory\[119\]\[2\] _01623_ _01624_ _01835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06229__A2 _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08474__I0 u_arbiter.i_wb_cpu_rdt\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07977__A2 _03626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[59\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08064_ u_arbiter.i_wb_cpu_rdt\[11\] _03669_ _03678_ u_arbiter.i_wb_cpu_dbus_dat\[11\]
+ _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05276_ u_cpu.rf_ram.memory\[76\]\[1\] u_cpu.rf_ram.memory\[77\]\[1\] u_cpu.rf_ram.memory\[78\]\[1\]
+ u_cpu.rf_ram.memory\[79\]\[1\] _01577_ _01549_ _01767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_135_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07015_ _02953_ _03081_ _03082_ _00415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07729__A2 _03458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06401__A2 _02718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08966_ _04343_ _01106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07917_ u_cpu.rf_ram.memory\[112\]\[0\] _03596_ _03597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08897_ u_cpu.rf_ram.memory\[95\]\[6\] _04299_ _04306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09351__A1 _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08154__A2 u_arbiter.i_wb_cpu_rdt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09723__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07848_ _03539_ _03558_ _03559_ _00772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_17_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05912__A1 _02311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07779_ u_cpu.rf_ram.memory\[35\]\[6\] _03510_ _03517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10700__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09518_ u_cpu.rf_ram.memory\[100\]\[5\] _04654_ _04660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10790_ _01219_ io_in[4] u_cpu.rf_ram.memory\[59\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09873__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09449_ u_cpu.rf_ram.memory\[25\]\[6\] _04615_ _04622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10850__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09406__A2 _04595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07417__A1 _03161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07968__A2 _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05979__A1 _01372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06640__A2 _02864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10224_ _00670_ io_in[4] u_cpu.rf_ram.memory\[124\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10155_ _00601_ io_in[4] u_cpu.rf_ram.memory\[131\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08868__I _02496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10230__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10086_ _00532_ io_in[4] u_cpu.rf_ram.memory\[138\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09342__A1 _02475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08145__A2 _03742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10380__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05903__A1 _02332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05903__B2 _01409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08817__B _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08309__S _01436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10988_ _10988_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_43_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07656__A1 _03343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07959__A2 _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05130_ _01589_ _01621_ _01622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05061_ _01397_ _01553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06631__A2 _02864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08908__A1 _04286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09746__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08820_ u_cpu.cpu.immdec.imm11_7\[3\] _03798_ _04253_ _04254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_140_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06395__A1 _02492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08751_ _02581_ u_cpu.rf_ram.memory\[3\]\[1\] _04208_ _04210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05963_ _01403_ _02422_ _02430_ _00014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10723__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08136__A2 _03731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09333__A1 _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07702_ u_cpu.rf_ram.memory\[91\]\[4\] _03465_ _03470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04914_ _01435_ _01436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08682_ u_cpu.cpu.ctrl.o_ibus_adr\[12\] _04155_ _04157_ u_cpu.cpu.ctrl.o_ibus_adr\[13\]
+ _04170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05894_ u_cpu.cpu.state.o_cnt_r\[1\] _02376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09896__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07633_ u_cpu.rf_ram.memory\[38\]\[7\] _03422_ _03430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04845_ _01369_ _01370_ u_cpu.cpu.bne_or_bge _01371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_54_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07564_ _03391_ _03392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10873__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05370__A2 _01859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09303_ _04482_ _04526_ _04533_ _01253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06515_ _02754_ _02791_ _02799_ _00198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07495_ u_cpu.rf_ram.memory\[22\]\[3\] _03345_ _03352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06446_ u_cpu.rf_ram.memory\[50\]\[6\] _02740_ _02753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09234_ _04484_ _04487_ _04495_ _01222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10103__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09165_ u_cpu.rf_ram.memory\[108\]\[4\] _04449_ _04454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06377_ _02492_ _02708_ _02711_ _00148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08116_ _03723_ _03678_ _03683_ _03725_ _03726_ _00873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__04881__A1 u_cpu.cpu.immdec.imm19_12_20\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05328_ _01422_ _01808_ _01817_ _01818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_134_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09096_ _04292_ _04409_ _04415_ _01164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08072__A1 u_arbiter.i_wb_cpu_rdt\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08072__B2 u_arbiter.i_wb_cpu_dbus_dat\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08047_ _03680_ _03681_ _00849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05259_ _01743_ _01745_ _01747_ _01749_ _01607_ _01750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__06622__A2 _02854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10253__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08375__A2 u_arbiter.i_wb_cpu_rdt\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09998_ _00005_ io_in[4] u_cpu.rf_ram.rdata\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08949_ u_arbiter.i_wb_cpu_rdt\[19\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[3\]
+ _04331_ _04335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08127__A2 _03731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09324__A1 _02475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05326__B _01626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10911_ _01340_ io_in[4] u_cpu.rf_ram.memory\[100\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10842_ _01271_ io_in[4] u_cpu.rf_ram.memory\[88\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07638__A1 _03343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10773_ _01202_ io_in[4] u_cpu.rf_ram.memory\[69\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09619__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05996__B _02332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06861__A2 _02992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09769__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07810__A1 _03351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05416__A3 _01904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06613__A2 _02854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10746__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09563__A1 _02321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10207_ _00653_ io_in[4] u_cpu.rf_ram.memory\[126\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06377__A1 _02492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10138_ _00584_ io_in[4] u_cpu.rf_ram.memory\[133\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09315__A1 _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08118__A2 _02781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10069_ _00515_ io_in[4] u_cpu.rf_ram.memory\[143\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10896__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10126__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06300_ u_cpu.rf_ram.memory\[45\]\[3\] _02662_ _02666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07280_ u_cpu.rf_ram.memory\[138\]\[5\] _03225_ _03231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06301__A1 _02497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05104__A2 _01595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06231_ _02522_ _02623_ _02624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10276__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04863__A1 u_cpu.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06162_ _02573_ u_cpu.rf_ram.memory\[1\]\[0\] _02578_ _02579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05113_ _01416_ _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06604__A2 _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07801__A1 _02524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06093_ _02507_ _02530_ _02536_ _00039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05044_ u_cpu.cpu.ctrl.o_ibus_adr\[31\] _01536_ _01537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09921_ _00375_ io_in[4] u_cpu.rf_ram.memory\[58\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08357__A2 _03931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09852_ _00306_ io_in[4] u_cpu.rf_ram.memory\[65\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06368__A1 _02517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08803_ _02312_ _04237_ _04238_ _04010_ _01048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_86_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09783_ _00237_ io_in[4] u_cpu.rf_ram.memory\[139\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06995_ _03070_ _03071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09306__A1 _02727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08109__A2 _03653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08734_ u_cpu.rf_ram.memory\[109\]\[1\] _04199_ _04201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05946_ _02320_ _02420_ _02421_ _00019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_96_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05591__A2 _02073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07868__A1 _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05877_ _02358_ _02308_ _02325_ _02359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_08665_ _04161_ _00987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_54_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07616_ _03359_ _03412_ _03420_ _00678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06540__A1 _02742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08596_ _04120_ _00959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_41_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07547_ u_cpu.rf_ram.memory\[126\]\[0\] _03382_ _03383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10619__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07478_ _03340_ _00620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07096__A2 _03119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09217_ _02684_ _02706_ _04486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06843__A2 _02982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06429_ _02738_ _02740_ _02741_ _00170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_6_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09911__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08192__B _03791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08045__A1 u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09148_ _04290_ _04439_ _04444_ _01187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10769__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09079_ u_cpu.rf_ram.memory\[79\]\[6\] _04399_ _04406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11110_ io_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_123_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11041_ _11041_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__09545__A1 _04468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07020__A2 _03081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05582__A2 _02064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10149__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06906__I0 _02573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08367__B _03763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08520__A2 _03798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06531__A1 _02752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10825_ _01254_ io_in[4] u_cpu.rf_ram.memory\[86\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08808__B1 _03779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05503__C _01628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10299__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08284__A1 _03756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07087__A2 _03119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10756_ _01185_ io_in[4] u_cpu.rf_ram.memory\[83\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08284__B2 _03867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09591__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10687_ _01116_ io_in[4] u_cpu.rf_ram.memory\[101\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__04845__A1 _01369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05193__S1 _01681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07497__I _02501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04914__I _01435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08036__A1 _03668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06598__A1 _02744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07011__A2 _03071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05800_ u_cpu.rf_ram.memory\[68\]\[7\] u_cpu.rf_ram.memory\[69\]\[7\] u_cpu.rf_ram.memory\[70\]\[7\]
+ u_cpu.rf_ram.memory\[71\]\[7\] _01555_ _01652_ _02285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_49_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06780_ _02746_ _02944_ _02948_ _00314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_48_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05573__A2 _02055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06770__A1 _02754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05731_ _01406_ _02167_ _02216_ _00006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_82_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08511__A2 _04070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08450_ _03993_ _04016_ _04017_ _03855_ _00916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05662_ u_cpu.rf_ram.memory\[52\]\[6\] u_cpu.rf_ram.memory\[53\]\[6\] u_cpu.rf_ram.memory\[54\]\[6\]
+ u_cpu.rf_ram.memory\[55\]\[6\] _01590_ _01591_ _02148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_91_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07401_ _03163_ _03295_ _03298_ _00585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08381_ _03946_ _03953_ _03955_ _00909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05593_ _01539_ _02051_ _02060_ _02079_ _02080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_108_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09934__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07332_ u_cpu.rf_ram.memory\[49\]\[4\] _03255_ _03260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08275__A1 _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08275__B2 _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07263_ _03221_ _00524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10911__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06825__A2 _02972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06214_ u_cpu.rf_ram.memory\[80\]\[0\] _02614_ _02615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09002_ _04288_ _04359_ _04363_ _01122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08027__A1 u_arbiter.i_wb_cpu_dbus_dat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07194_ _03171_ _03176_ _03183_ _00493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06145_ u_cpu.rf_ram.memory\[20\]\[3\] _02563_ _02567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06076_ u_cpu.cpu.immdec.imm11_7\[4\] _02525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07250__A2 _03206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09527__A1 _04468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05027_ u_cpu.cpu.ctrl.o_ibus_adr\[27\] _01523_ _01524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09904_ _00358_ io_in[4] u_cpu.rf_ram.memory\[60\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07002__A2 _03071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09835_ _00289_ io_in[4] u_cpu.rf_ram.memory\[67\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05013__A1 u_arbiter.i_wb_cpu_dbus_adr\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09766_ _00220_ io_in[4] u_cpu.rf_ram.memory\[119\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06687__S _02894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06978_ u_cpu.rf_ram.memory\[55\]\[0\] _03061_ _03062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08717_ _04188_ _01012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_26_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05929_ _01374_ _02373_ _02409_ _01386_ _02410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09697_ _00151_ io_in[4] u_cpu.rf_ram.memory\[43\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10441__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08648_ u_cpu.rf_ram.memory\[30\]\[5\] _04145_ _04151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06513__A1 _02752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08579_ _04111_ _00951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10610_ _01039_ io_in[4] u_cpu.rf_ram.memory\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08266__A1 _03761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10591__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10541_ _00022_ io_in[4] u_cpu.cpu.bufreg.c_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08018__A1 u_arbiter.i_wb_cpu_dbus_dat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10472_ _00905_ io_in[4] u_cpu.cpu.immdec.imm24_20\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09238__S _04496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08142__S _01434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05993__C _02448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07241__A2 _03206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05252__A1 _01398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09807__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11024_ _11024_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08741__A2 _04199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05555__A2 _01993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06752__A1 _02754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09957__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[63\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10934__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10808_ _01237_ io_in[4] u_cpu.rf_ram.memory\[85\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08257__A1 _03786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06807__A2 _02955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10739_ _01168_ io_in[4] u_cpu.rf_ram.memory\[106\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05166__S1 _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08009__A1 u_arbiter.i_wb_cpu_dbus_dat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05491__A1 _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07232__A2 _03196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10314__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05243__A1 _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09509__A1 _04468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07950_ _03555_ _03606_ _03614_ _00819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08980__A2 _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06991__A1 _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06901_ u_cpu.rf_ram.memory\[19\]\[6\] _03012_ _03019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07881_ _02577_ _02810_ _03577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[16\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08732__A2 _04199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09620_ _00074_ io_in[4] u_cpu.rf_ram.memory\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09391__B _01393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06832_ _02969_ _02972_ _02980_ _00334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10464__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05546__A2 _02033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09551_ _04476_ _04674_ _04678_ _01356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06763_ u_cpu.rf_ram.memory\[65\]\[4\] _02934_ _02939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08502_ _04060_ _04062_ _03980_ _04063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05714_ u_cpu.rf_ram.memory\[72\]\[6\] u_cpu.rf_ram.memory\[73\]\[6\] u_cpu.rf_ram.memory\[74\]\[6\]
+ u_cpu.rf_ram.memory\[75\]\[6\] _01610_ _01611_ _02200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09482_ _02593_ u_cpu.rf_ram.memory\[0\]\[5\] _04634_ _04640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06694_ _02900_ _00276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_24_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07299__A2 _03235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08433_ _03999_ _04000_ _04001_ _03755_ _04002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_52_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05645_ _01542_ _02130_ _02131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08248__A1 _03757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08364_ _03934_ _03938_ _03939_ _00908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05576_ u_cpu.rf_ram.memory\[48\]\[5\] u_cpu.rf_ram.memory\[49\]\[5\] u_cpu.rf_ram.memory\[50\]\[5\]
+ u_cpu.rf_ram.memory\[51\]\[5\] _01544_ _01548_ _02063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08799__A2 _04227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07315_ _03167_ _03245_ _03250_ _00547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08295_ u_cpu.rf_ram.memory\[114\]\[2\] _03879_ _03882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07246_ _03169_ _03206_ _03212_ _00516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05482__A1 _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07177_ u_cpu.rf_ram.memory\[72\]\[7\] _03159_ _03174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06128_ _02502_ _02551_ _02556_ _00054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07223__A2 _03196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08420__A1 _03987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05234__A1 _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06059_ _02460_ u_cpu.rf_ram_if.wdata0_r\[6\] _02509_ _02510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_78_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10807__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05318__C _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09818_ _00272_ io_in[4] u_cpu.rf_ram.memory\[6\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08723__A2 _01386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06734__A1 _02754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09749_ _00203_ io_in[4] u_cpu.rf_ram.memory\[17\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08487__A1 _04016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08239__A1 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10524_ _00957_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07462__A2 _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10337__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05473__A1 _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10455_ _00888_ io_in[4] u_cpu.cpu.branch_op vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07214__A2 _03186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08411__A1 _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10386_ _00819_ io_in[4] u_cpu.rf_ram.memory\[122\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05225__A1 _01594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[22\] u_arbiter.i_wb_cpu_rdt\[19\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[16\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__05509__B _01416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10487__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06973__A1 _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11007_ _11007_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__08714__A2 _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05528__A2 _02015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08478__A1 _03756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05430_ _01645_ _01918_ _01648_ _01919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05700__A2 _02176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05361_ _01553_ _01850_ _01565_ _01851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_105_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07886__S _03577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07100_ _02660_ _02832_ _03128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08080_ u_arbiter.i_wb_cpu_rdt\[17\] _03653_ _03654_ u_arbiter.i_wb_cpu_dbus_dat\[17\]
+ _03676_ u_arbiter.i_wb_cpu_dbus_dat\[18\] _03703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_05292_ u_cpu.rf_ram.memory\[8\]\[2\] u_cpu.rf_ram.memory\[9\]\[2\] u_cpu.rf_ram.memory\[10\]\[2\]
+ u_cpu.rf_ram.memory\[11\]\[2\] _01546_ _01550_ _01782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07453__A2 _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07031_ _03090_ _03091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05464__A1 _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08402__A1 _03973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07205__A2 _03186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05216__A1 _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08982_ _04286_ _04349_ _04352_ _01113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07933_ _02638_ _02821_ _03605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07864_ _03567_ _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06716__A1 _02754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09603_ _00057_ io_in[4] u_cpu.rf_ram.memory\[18\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06815_ _02684_ _02727_ _02971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07795_ u_cpu.rf_ram.memory\[34\]\[5\] _03520_ _03526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09534_ u_cpu.rf_ram.memory\[89\]\[4\] _04664_ _04669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06746_ _02748_ _02924_ _02929_ _00299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09130__A2 _04429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09465_ u_cpu.rf_ram.memory\[24\]\[5\] _04625_ _04631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06677_ u_cpu.rf_ram.memory\[75\]\[6\] _02884_ _02891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08416_ _03742_ _03751_ _03741_ _03986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05628_ u_cpu.rf_ram.memory\[76\]\[5\] u_cpu.rf_ram.memory\[77\]\[5\] u_cpu.rf_ram.memory\[78\]\[5\]
+ u_cpu.rf_ram.memory\[79\]\[5\] _01577_ _01549_ _02115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07692__A2 _02706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09396_ _03812_ _04592_ _01287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08347_ _03831_ _03790_ _03818_ _03819_ _03924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_138_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05559_ _01554_ _02045_ _01417_ _02046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09652__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08278_ _03801_ _03858_ _03868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07444__A2 _03315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08641__A1 _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05455__A1 _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07229_ u_cpu.rf_ram.memory\[70\]\[6\] _03196_ _03203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09197__A2 _04470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10240_ _00009_ io_in[4] u_cpu.rf_ram_if.rdata0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06205__S _02603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05207__A1 _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10171_ _00617_ io_in[4] u_cpu.rf_ram.memory\[12\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06955__A1 _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05066__S0 _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04887__C _01377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09121__A2 _04429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05999__B u_cpu.rf_ram_if.genblk1.wtrig0_r vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05369__S1 _01681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07683__A2 _03458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05694__A1 _01601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07435__A2 _03315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10507_ _00940_ io_in[4] u_cpu.rf_ram.memory\[31\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05997__A2 _02431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09188__A2 _04459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10438_ _00871_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08935__A2 _04322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10369_ _00802_ io_in[4] u_cpu.rf_ram.memory\[11\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04930_ u_arbiter.i_wb_cpu_dbus_adr\[4\] _01443_ _01450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09360__A2 _01386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04861_ _01379_ _01382_ _01386_ _01387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07371__A1 _03169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06600_ _02746_ _02844_ _02848_ _00234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07580_ _03359_ _03392_ _03400_ _00662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_19_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05921__A2 _02401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09112__A2 _04419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06531_ _02752_ _02801_ _02808_ _00205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10502__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07123__A1 _02957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09250_ _02599_ u_cpu.rf_ram.memory\[10\]\[7\] _04496_ _04504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09675__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06462_ _02593_ u_cpu.rf_ram.memory\[4\]\[5\] _02756_ _02762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07674__A2 u_cpu.cpu.state.o_cnt_r\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05685__A1 _01594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08201_ _02765_ u_arbiter.i_wb_cpu_rdt\[1\] _03799_ _03800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_33_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05413_ u_cpu.rf_ram.memory\[32\]\[3\] u_cpu.rf_ram.memory\[33\]\[3\] u_cpu.rf_ram.memory\[34\]\[3\]
+ u_cpu.rf_ram.memory\[35\]\[3\] _01623_ _01624_ _01902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09181_ u_cpu.rf_ram.memory\[69\]\[3\] _04459_ _04463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06393_ _02487_ _02718_ _02720_ _00155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08132_ u_cpu.rf_ram.memory\[113\]\[4\] _03731_ _03736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10652__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05344_ _01541_ _01833_ _01834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07426__A2 _03305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08474__I1 u_arbiter.i_wb_cpu_rdt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08063_ u_arbiter.i_wb_cpu_dbus_dat\[12\] _03683_ _03692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05275_ _01667_ _01765_ _01766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07014_ u_cpu.rf_ram.memory\[53\]\[0\] _03081_ _03082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09179__A2 _04459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08926__A2 _04322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[9\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06937__A1 _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05296__S0 _01546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08965_ u_arbiter.i_wb_cpu_rdt\[27\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[11\]
+ _04331_ _04343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07916_ _03595_ _03596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10032__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08896_ _04292_ _04299_ _04305_ _01074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__04963__A3 _01462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09351__A2 _04556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07847_ u_cpu.rf_ram.memory\[118\]\[0\] _03558_ _03559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06695__S _02894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07778_ _03355_ _03510_ _03516_ _00745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10182__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09103__A2 _04419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09517_ _04478_ _04654_ _04659_ _01341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06729_ u_cpu.rf_ram.memory\[67\]\[5\] _02914_ _02920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08162__I0 u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09448_ _04480_ _04615_ _04621_ _01310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07665__A2 _03442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05676__A1 _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09379_ u_cpu.cpu.genblk3.csr.mcause31 _04580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_32_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08415__S _01437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07417__A2 _03305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05428__A1 _01398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05979__A2 _02394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08917__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10223_ _00669_ io_in[4] u_cpu.rf_ram.memory\[124\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09246__S _04496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05287__S0 _01687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10154_ _00600_ io_in[4] u_cpu.rf_ram.memory\[131\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10085_ _00531_ io_in[4] u_cpu.rf_ram.memory\[138\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09342__A2 _02810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08145__A3 _03743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10525__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07353__A1 _03169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09698__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05903__A2 u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10987_ _10987_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_90_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07105__A1 _02957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05522__B _01654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10675__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07656__A2 _03442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05667__A1 _01636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07408__A2 _03295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05419__A1 _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05060_ _01542_ _01551_ _01552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08908__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10055__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07592__A1 _03353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06395__A2 _02718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08750_ _04209_ _01024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05962_ u_cpu.rf_ram_if.rdata0\[7\] _01403_ _02430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07701_ _03351_ _03465_ _03469_ _00714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09333__A2 _04546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04913_ _01434_ _01435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08681_ _04169_ _00995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_94_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06147__A2 _02563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05893_ _02354_ _02374_ _01373_ _02363_ _02375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_65_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07632_ _03357_ _03422_ _03429_ _00685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_4_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04844_ u_cpu.cpu.decode.co_mem_word _01370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05450__S0 _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07563_ _02660_ _02821_ _03391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08144__I0 u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09302_ u_cpu.rf_ram.memory\[86\]\[6\] _04526_ _04533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06514_ u_cpu.rf_ram.memory\[16\]\[7\] _02791_ _02799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08844__A1 _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07647__A2 _03432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[26\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07494_ _02496_ _03351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05658__A1 _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09233_ u_cpu.rf_ram.memory\[59\]\[7\] _04487_ _04495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06445_ _02511_ _02752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09164_ _04288_ _04449_ _04453_ _01194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06376_ u_cpu.rf_ram.memory\[43\]\[2\] _02708_ _02711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08235__S _01435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06458__I0 _02587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08115_ u_arbiter.i_wb_cpu_rdt\[29\] _02781_ _03726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__04881__A2 u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05327_ _01810_ _01812_ _01814_ _01816_ _01628_ _01817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_09095_ u_cpu.rf_ram.memory\[105\]\[5\] _04409_ _04415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08072__A2 _03653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06083__A1 _02482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08046_ u_arbiter.i_wb_cpu_dbus_dat\[5\] _03654_ _03676_ _02779_ _03681_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05258_ _01614_ _01748_ _01654_ _01749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05830__A1 _01372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05189_ _01668_ _01681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09997_ _00004_ io_in[4] u_cpu.rf_ram.rdata\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10548__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06386__A2 _02708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08948_ _04334_ _01097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09840__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09324__A2 _02602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08879_ _04294_ _04282_ _04295_ _01067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07335__A1 _03169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10910_ _01339_ io_in[4] u_cpu.rf_ram.memory\[100\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10698__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05441__S0 _01590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05897__A1 _02338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10841_ _01270_ io_in[4] u_cpu.rf_ram.memory\[87\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09088__A1 _04284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09990__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05342__B _01648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07638__A2 _03432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10772_ _01201_ io_in[4] u_cpu.rf_ram.memory\[69\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05649__A1 _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06697__I0 _02599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08048__C1 _03676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10078__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08063__A2 _03683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07810__A2 _03530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10206_ _00652_ io_in[4] u_cpu.rf_ram.memory\[126\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09563__A2 _02320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07574__A1 _03353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06377__A2 _02708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10137_ _00583_ io_in[4] u_cpu.rf_ram.memory\[133\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09315__A2 _04536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10068_ _00514_ io_in[4] u_cpu.rf_ram.memory\[143\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06129__A2 _02551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07877__A2 _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[49\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05888__A1 u_cpu.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07629__A2 _03422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08826__A1 _03755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06301__A2 _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06230_ _01386_ _02462_ _02623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_54_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04863__A2 _01388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09713__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06161_ _02539_ _02577_ _02578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08054__A2 _03683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07894__S _03577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06065__A1 _02460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05499__S0 _01619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05112_ u_cpu.rf_ram.memory\[56\]\[0\] u_cpu.rf_ram.memory\[57\]\[0\] u_cpu.rf_ram.memory\[58\]\[0\]
+ u_cpu.rf_ram.memory\[59\]\[0\] _01602_ _01603_ _01604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_06092_ u_cpu.rf_ram.memory\[21\]\[5\] _02530_ _02536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07801__A2 _02821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05043_ _01535_ _01532_ _01536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09920_ _00374_ io_in[4] u_cpu.rf_ram.memory\[5\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05812__A1 _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09863__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09554__A2 _04674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09851_ _00305_ io_in[4] u_cpu.rf_ram.memory\[65\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06368__A2 _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08802_ u_cpu.cpu.immdec.imm11_7\[1\] _03797_ _04237_ _04238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09782_ _00236_ io_in[4] u_cpu.rf_ram.memory\[139\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06994_ _02684_ _02893_ _03070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10840__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05040__A2 _01457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08733_ _03539_ _04199_ _04200_ _01016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09306__A2 _04197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05671__S0 _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05945_ _02320_ u_cpu.rf_ram_if.rdata1\[5\] _02421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07317__A1 _03169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08664_ u_cpu.cpu.ctrl.o_ibus_adr\[3\] _04155_ _04157_ u_cpu.cpu.ctrl.o_ibus_adr\[4\]
+ _04161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_26_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07868__A2 _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05876_ _02309_ u_cpu.cpu.alu.add_cy_r _02358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_26_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07615_ u_cpu.rf_ram.memory\[123\]\[7\] _03412_ _03420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08595_ u_arbiter.i_wb_cpu_dbus_adr\[18\] u_arbiter.i_wb_cpu_dbus_adr\[17\] _04115_
+ _04120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06540__A2 _02812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07546_ _03381_ _03382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08817__A1 _03810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08293__A2 _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07477_ _02593_ u_cpu.rf_ram.memory\[12\]\[5\] _03334_ _03340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10220__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09216_ _04484_ _04470_ _04485_ _01214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06428_ u_cpu.rf_ram.memory\[50\]\[0\] _02740_ _02741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09147_ u_cpu.rf_ram.memory\[83\]\[4\] _04439_ _04444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06359_ u_cpu.rf_ram.memory\[41\]\[3\] _02697_ _02701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08045__A2 _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09078_ _04292_ _04399_ _04405_ _01156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10370__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05803__A1 _01609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08029_ u_arbiter.i_wb_cpu_rdt\[2\] _02781_ _03666_ _03667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11040_ _11040_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__09545__A2 _04674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07556__A1 _03353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06359__A2 _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05337__B _01626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05662__S0 _01590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07859__A2 _03558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06531__A2 _02801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10824_ _01253_ io_in[4] u_cpu.rf_ram.memory\[86\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08808__A1 _03761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08808__B2 _03788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10755_ _01184_ io_in[4] u_cpu.rf_ram.memory\[83\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09736__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08284__A2 _03778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06295__A1 _02482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10686_ _01115_ io_in[4] u_cpu.rf_ram.memory\[101\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10713__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[52\] u_scanchain_local.module_data_in\[51\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[14\] u_scanchain_local.clk u_scanchain_local.module_data_in\[52\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__04845__A2 _01370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08036__A2 _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06047__A1 _02460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09886__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08603__S _04115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06598__A2 _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10863__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09536__A2 _04664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05653__S0 _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06770__A2 _02934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05730_ _02206_ _02215_ _02216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05661_ _02140_ _02142_ _02144_ _02146_ _01426_ _02147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_90_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06522__A2 _02801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10243__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07400_ u_cpu.rf_ram.memory\[133\]\[2\] _03295_ _03298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08380_ u_cpu.cpu.immdec.imm30_25\[0\] _03954_ _03955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05592_ _01422_ _02069_ _02078_ _02079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_07331_ _03165_ _03255_ _03259_ _00554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08275__A2 _03856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06286__A1 _02507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07262_ _02593_ u_cpu.rf_ram.memory\[14\]\[5\] _03215_ _03221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10393__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09001_ u_cpu.rf_ram.memory\[102\]\[3\] _04359_ _04363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06213_ _02613_ _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07193_ u_cpu.rf_ram.memory\[73\]\[6\] _03176_ _03183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09224__A1 _04474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06144_ _02492_ _02563_ _02566_ _00060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07786__A1 _03343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06589__A2 _02834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06075_ _02521_ _02523_ _02524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05797__B1 _02279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09527__A2 _04664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05026_ u_cpu.cpu.ctrl.o_ibus_adr\[26\] u_cpu.cpu.ctrl.o_ibus_adr\[25\] u_cpu.cpu.ctrl.o_ibus_adr\[24\]
+ _01513_ _01523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_09903_ _00357_ io_in[4] u_cpu.rf_ram.memory\[60\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07538__A1 _03353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05157__B _01648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09834_ _00288_ io_in[4] u_cpu.rf_ram.memory\[67\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09609__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05013__A2 _01442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05644__S0 _01546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09765_ _00219_ io_in[4] u_cpu.rf_ram.memory\[119\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06977_ _03060_ _03061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_58_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06761__A2 _02934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08716_ u_cpu.cpu.ctrl.o_ibus_adr\[28\] _04173_ _04175_ u_cpu.cpu.ctrl.o_ibus_adr\[29\]
+ _04188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_100_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05928_ _01374_ _02406_ _02409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09696_ _00150_ io_in[4] u_cpu.rf_ram.memory\[43\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08647_ _03549_ _04145_ _04150_ _00980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09759__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05859_ _02311_ u_cpu.cpu.genblk3.csr.mcause31 _02338_ _02342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07710__A1 _02475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06513__A2 _02791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08578_ u_arbiter.i_wb_cpu_dbus_adr\[10\] u_arbiter.i_wb_cpu_dbus_adr\[9\] _02445_
+ _04111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07529_ u_cpu.rf_ram.memory\[127\]\[0\] _03372_ _03373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10736__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08266__A2 _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05620__B _01654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10540_ _00973_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08018__A2 u_arbiter.i_wb_cpu_dbus_dat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10471_ _00904_ io_in[4] u_cpu.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06029__A1 _02460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10886__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05252__A2 _01742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09518__A2 _04654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10116__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11023_ _11023_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_110_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05067__B _01417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05635__S0 _01680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06752__A2 _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10266__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05514__C _01628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07701__A1 _03351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06504__A2 _02791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10807_ _01236_ io_in[4] u_cpu.rf_ram.memory\[85\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08257__A2 _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06268__A1 _02507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10738_ _01167_ io_in[4] u_cpu.rf_ram.memory\[106\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08009__A2 _02774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10669_ _01098_ io_in[4] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07068__I0 _02581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05491__A2 _01978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07768__A1 _03343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05243__A2 _01733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09509__A2 _04654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06991__A2 _03061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06900_ _02965_ _03012_ _03018_ _00364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07880_ _03555_ _03568_ _03576_ _00787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10609__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08193__A1 _03752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06831_ u_cpu.rf_ram.memory\[63\]\[7\] _02972_ _02980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05626__S0 _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08288__B _03877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06743__A2 _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07940__A1 _03545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09901__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09550_ u_cpu.rf_ram.memory\[23\]\[3\] _04674_ _04678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06762_ _02746_ _02934_ _02938_ _00306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08501_ _03742_ _03897_ _04061_ _03791_ _04062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05713_ _01553_ _02198_ _01565_ _02199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_58_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10759__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09481_ _04639_ _01325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06693_ _02593_ u_cpu.rf_ram.memory\[6\]\[5\] _02894_ _02900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08496__A2 _04016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08432_ _03749_ _03831_ _03770_ _04001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_23_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05644_ u_cpu.rf_ram.memory\[8\]\[6\] u_cpu.rf_ram.memory\[9\]\[6\] u_cpu.rf_ram.memory\[10\]\[6\]
+ u_cpu.rf_ram.memory\[11\]\[6\] _01546_ _01550_ _02130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_63_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08363_ u_cpu.cpu.immdec.imm24_20\[4\] _03916_ _03919_ u_cpu.cpu.immdec.imm30_25\[0\]
+ _03935_ _03816_ _03939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__08248__A2 _03759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05575_ _01589_ _02061_ _02062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05440__B _01648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07314_ u_cpu.rf_ram.memory\[137\]\[4\] _03245_ _03250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08294_ _03543_ _03879_ _03881_ _00896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07245_ u_cpu.rf_ram.memory\[143\]\[5\] _03206_ _03212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07059__I0 _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10139__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07176_ _02516_ _03173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_106_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06127_ u_cpu.rf_ram.memory\[18\]\[4\] _02551_ _02556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05234__A2 _01724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08042__I _03654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06058_ _02478_ u_cpu.rf_ram_if.wdata1_r\[6\] _02509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_8_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08708__B1 _04175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06982__A2 _03061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10289__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05009_ _01443_ _01508_ _01509_ _01510_ u_arbiter.o_wb_cpu_adr\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_143_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08184__A1 _01435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05617__S0 _01590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09817_ _00271_ io_in[4] u_cpu.rf_ram.memory\[6\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09581__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06734__A2 _02914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09748_ _00202_ io_in[4] u_cpu.rf_ram.memory\[17\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09679_ _00133_ io_in[4] u_cpu.rf_ram.memory\[51\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06498__A1 _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07998__A1 _03549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10523_ _00956_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05473__A2 _01960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06670__A1 _02744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10454_ _00887_ io_in[4] u_arbiter.i_wb_cpu_dbus_we vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10385_ _00818_ io_in[4] u_cpu.rf_ram.memory\[122\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06422__A1 _02512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05225__A2 _01715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06973__A2 _03051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09924__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[15\] u_arbiter.i_wb_cpu_rdt\[12\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[9\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_46_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11006_ _11006_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_93_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10901__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07922__A1 _03545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06725__A2 _02914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.input_buf_clk io_in[0] u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_92_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05700__A3 _02185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05360_ u_cpu.rf_ram.memory\[68\]\[2\] u_cpu.rf_ram.memory\[69\]\[2\] u_cpu.rf_ram.memory\[70\]\[2\]
+ u_cpu.rf_ram.memory\[71\]\[2\] _01555_ _01652_ _01850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_119_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05291_ _01406_ _01732_ _01781_ _00001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08650__A2 _04145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07030_ _02561_ _02684_ _03090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05464__A2 _01952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08402__A2 _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10431__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05216__A2 _01706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08981_ u_cpu.rf_ram.memory\[101\]\[2\] _04349_ _04352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06964__A2 _03051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07932_ _03555_ _03596_ _03604_ _00811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04975__A1 u_cpu.cpu.ctrl.o_ibus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08166__A1 _01435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07863_ _02695_ _02821_ _03567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10581__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06716__A2 _02904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08961__I0 u_arbiter.i_wb_cpu_rdt\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06814_ _02969_ _02955_ _02970_ _00326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09602_ _00056_ io_in[4] u_cpu.rf_ram.memory\[18\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07794_ _03353_ _03520_ _03525_ _00752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09533_ _04476_ _04664_ _04668_ _01348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06745_ u_cpu.rf_ram.memory\[66\]\[4\] _02924_ _02929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09464_ _04478_ _04625_ _04630_ _01317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06676_ _02750_ _02884_ _02890_ _00268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08415_ u_arbiter.i_wb_cpu_rdt\[30\] u_arbiter.i_wb_cpu_rdt\[14\] _01437_ _03985_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05627_ _01667_ _02113_ _02114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05152__A1 _01398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09395_ u_cpu.cpu.ctrl.i_iscomp _03798_ _04592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08346_ u_arbiter.i_wb_cpu_rdt\[23\] u_arbiter.i_wb_cpu_rdt\[7\] _01436_ _03923_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_138_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05558_ u_cpu.rf_ram.memory\[12\]\[5\] u_cpu.rf_ram.memory\[13\]\[5\] u_cpu.rf_ram.memory\[14\]\[5\]
+ u_cpu.rf_ram.memory\[15\]\[5\] _01556_ _01557_ _02045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_138_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08277_ u_arbiter.i_wb_cpu_rdt\[22\] u_arbiter.i_wb_cpu_rdt\[6\] _01436_ _03867_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05489_ _01594_ _01976_ _01564_ _01977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08641__A2 _04145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08481__B _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05455__A2 _01934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06652__A1 _02744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07228_ _03169_ _03196_ _03202_ _00508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09947__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07159_ u_cpu.rf_ram.memory\[72\]\[1\] _03159_ _03162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05207__A2 _01697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10170_ _00616_ io_in[4] u_cpu.rf_ram.memory\[12\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_u_scanchain_local.scan_flop\[62\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10924__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06955__A2 _03041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06707__A2 _02904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05066__S1 _01557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07380__A2 _03285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07132__A2 _03139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10304__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05143__A1 _01594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[15\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08632__A2 _02448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10454__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10506_ _00939_ io_in[4] u_cpu.rf_ram.memory\[31\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10437_ _00870_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08396__A1 _02765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07199__A2 _03186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10368_ _00801_ io_in[4] u_cpu.rf_ram.memory\[11\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08611__S _04115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05239__C _01628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06946__A2 _03041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10299_ _00732_ io_in[4] u_cpu.rf_ram.memory\[92\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08943__I0 u_arbiter.i_wb_cpu_rdt\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[7\]_SI u_arbiter.i_wb_cpu_dbus_dat\[1\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04860_ _01378_ _01383_ _01384_ _01385_ _01386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_20_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07371__A2 _03275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06530_ u_cpu.rf_ram.memory\[17\]\[6\] _02801_ _02808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08320__A1 _03741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07123__A2 _03139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06461_ _02761_ _00182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06182__I0 _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08200_ _01436_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\] _03799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05412_ _01589_ _01900_ _01901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05685__A2 _02170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06882__A1 _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09180_ _04286_ _04459_ _04462_ _01201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06392_ u_cpu.rf_ram.memory\[48\]\[1\] _02718_ _02720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08131_ _03547_ _03731_ _03735_ _00879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_18_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05343_ u_cpu.rf_ram.memory\[112\]\[2\] u_cpu.rf_ram.memory\[113\]\[2\] u_cpu.rf_ram.memory\[114\]\[2\]
+ u_cpu.rf_ram.memory\[115\]\[2\] _01619_ _01591_ _01833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_18_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08623__A2 _02445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06634__A1 _02744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08062_ _03690_ _03691_ _00854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05274_ u_cpu.rf_ram.memory\[72\]\[1\] u_cpu.rf_ram.memory\[73\]\[1\] u_cpu.rf_ram.memory\[74\]\[1\]
+ u_cpu.rf_ram.memory\[75\]\[1\] _01571_ _01668_ _01765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_134_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10947__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07013_ _03080_ _03081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08387__A1 _03773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05149__C _01628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06937__A2 _03031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05296__S1 _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08964_ _04342_ _01105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08139__A1 _03555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07137__S _03148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07915_ _02612_ _02821_ _03595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08895_ u_cpu.rf_ram.memory\[95\]\[5\] _04299_ _04305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07846_ _03557_ _03558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07362__A2 _03275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10327__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07777_ u_cpu.rf_ram.memory\[35\]\[5\] _03510_ _03516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04989_ u_cpu.cpu.ctrl.o_ibus_adr\[18\] u_cpu.cpu.ctrl.o_ibus_adr\[17\] u_cpu.cpu.ctrl.o_ibus_adr\[16\]
+ _01488_ _01495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_37_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08476__B _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09516_ u_cpu.rf_ram.memory\[100\]\[4\] _04654_ _04659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06728_ _02748_ _02914_ _02919_ _00291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08311__A1 _03785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07114__A2 _03129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09447_ u_cpu.rf_ram.memory\[25\]\[5\] _04615_ _04621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06659_ u_cpu.rf_ram.memory\[76\]\[6\] _02874_ _02881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10477__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09378_ _04578_ _04568_ _04579_ _02349_ _01282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_36_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08329_ _03767_ _03890_ _03769_ _03888_ _03826_ _03744_ _03910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XFILLER_36_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08075__B1 _03678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05428__A2 _01916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10222_ _00668_ io_in[4] u_cpu.rf_ram.memory\[124\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06928__A2 _03031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05287__S1 _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10153_ _00599_ io_in[4] u_cpu.rf_ram.memory\[131\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10084_ _00530_ io_in[4] u_cpu.rf_ram.memory\[138\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[8\] u_arbiter.i_wb_cpu_rdt\[5\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[2\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_43_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08145__A4 _03744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07353__A2 _03265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10986_ _10986_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__08302__A1 _03551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07105__A2 _03129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05116__A1 _01593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08853__A2 _04271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05667__A2 _02152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06864__A1 _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05419__A2 _01907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06616__A1 _02744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06092__A2 _02530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08369__A1 _03773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07041__A1 _02963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07592__A2 _03402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08140__I _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05961_ _01403_ _02420_ _02429_ _00013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07700_ u_cpu.rf_ram.memory\[91\]\[3\] _03465_ _03469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04912_ u_cpu.cpu.genblk1.align.ctrl_misal _01434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08680_ u_cpu.cpu.ctrl.o_ibus_adr\[11\] _04155_ _04157_ u_cpu.cpu.ctrl.o_ibus_adr\[12\]
+ _04169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_94_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05892_ _01370_ _02357_ _02360_ _02373_ _02374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_65_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09642__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08541__A1 _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07344__A2 _03265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07631_ u_cpu.rf_ram.memory\[38\]\[6\] _03422_ _03429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04843_ u_cpu.cpu.csr_d_sel _01369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07562_ _03359_ _03382_ _03390_ _00654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05713__B _01565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05450__S1 _01668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09097__A2 _04409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09301_ _04480_ _04526_ _04532_ _01252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_59_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06513_ _02752_ _02791_ _02798_ _00197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09792__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07493_ _03349_ _03345_ _03350_ _00625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08844__A2 _04271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09232_ _04482_ _04487_ _04494_ _01221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06444_ _02750_ _02740_ _02751_ _00175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05658__A2 _02143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09163_ u_cpu.rf_ram.memory\[108\]\[3\] _04449_ _04453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06375_ _02487_ _02708_ _02710_ _00147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08114_ u_arbiter.i_wb_cpu_dbus_dat\[30\] _03725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05326_ _01541_ _01815_ _01626_ _01816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_108_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09094_ _04290_ _04409_ _04414_ _01163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08045_ u_arbiter.i_wb_cpu_rdt\[5\] _03669_ _03680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06083__A2 _02530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05257_ u_cpu.rf_ram.memory\[116\]\[1\] u_cpu.rf_ram.memory\[117\]\[1\] u_cpu.rf_ram.memory\[118\]\[1\]
+ u_cpu.rf_ram.memory\[119\]\[1\] _01623_ _01624_ _01748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_122_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05830__A2 u_cpu.cpu.decode.opcode\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09021__A2 _04369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05188_ _01571_ _01680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_1_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09996_ _00003_ io_in[4] u_cpu.rf_ram.rdata\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07583__A2 _03402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08050__I _03676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08947_ u_arbiter.i_wb_cpu_rdt\[18\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[2\]
+ _04331_ _04334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08878_ u_cpu.rf_ram.memory\[94\]\[6\] _04282_ _04295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07335__A2 _03255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07829_ _03545_ _03541_ _03546_ _00766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05346__A1 _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10840_ _01269_ io_in[4] u_cpu.rf_ram.memory\[87\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05441__S1 _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09088__A2 _04409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07099__A1 _02969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10771_ _01200_ io_in[4] u_cpu.rf_ram.memory\[69\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08835__A2 _03809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05649__A2 _02134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06846__A1 _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07894__I0 _02596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08048__B1 _03654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05849__I _01370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09260__A2 _04506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07271__A1 _03157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10205_ _00651_ io_in[4] u_cpu.rf_ram.memory\[126\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07023__A1 _02963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09665__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07574__A2 _03392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10136_ _00582_ io_in[4] u_cpu.rf_ram.memory\[134\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10067_ _00513_ io_in[4] u_cpu.rf_ram.memory\[143\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10642__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08523__A1 _02311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07326__A2 _03255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05337__A1 _01601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09079__A2 _04399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10792__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10969_ _10969_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__08826__A2 _03786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[8\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10022__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06160_ _02576_ _02577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05111_ _01547_ _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06065__A2 u_cpu.cpu.o_wdata0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05499__S1 _01620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06091_ _02502_ _02530_ _02535_ _00038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05042_ u_cpu.cpu.ctrl.o_ibus_adr\[30\] _01535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_144_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09003__A2 _04359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10172__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05708__B _01654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09850_ _00304_ io_in[4] u_cpu.rf_ram.memory\[65\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07565__A2 _03392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08801_ _02768_ _04236_ _04237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_140_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05120__S0 _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06993_ _02969_ _03061_ _03069_ _00406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09781_ _00235_ io_in[4] u_cpu.rf_ram.memory\[139\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08732_ u_cpu.rf_ram.memory\[109\]\[0\] _04199_ _04200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05944_ _02321_ u_cpu.rf_ram.rdata\[5\] _02420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05671__S1 _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08514__A1 _03797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07317__A2 _03245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08663_ _04160_ _00986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_22_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05328__A1 _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05875_ _01369_ _02355_ _02356_ _02357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_81_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07614_ _03357_ _03412_ _03419_ _00677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08594_ _04119_ _00958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07545_ _02625_ _02821_ _03381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06828__A1 _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07476_ _03339_ _00619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09490__A2 _04644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09215_ u_cpu.rf_ram.memory\[84\]\[7\] _04470_ _04485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06427_ _02739_ _02740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05500__A1 _01589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09146_ _04288_ _04439_ _04443_ _01186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06358_ _02492_ _02697_ _02700_ _00140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10515__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06056__A2 _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05309_ _01792_ _01794_ _01796_ _01798_ _01426_ _01799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_09077_ u_cpu.rf_ram.memory\[79\]\[5\] _04399_ _04405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06289_ u_cpu.rf_ram.memory\[46\]\[7\] _02651_ _02659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09688__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08028_ _03662_ _03664_ _02781_ _03665_ _03666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__05803__A2 _02287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07005__A1 _02963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10665__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07556__A2 _03382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09979_ _00433_ io_in[4] u_cpu.rf_ram.memory\[9\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05662__S1 _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07308__A2 _03245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10823_ _01252_ io_in[4] u_cpu.rf_ram.memory\[86\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08808__A2 _03778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10045__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10754_ _01183_ io_in[4] u_cpu.rf_ram.memory\[83\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08156__S _01435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06295__A2 _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10685_ _01114_ io_in[4] u_cpu.rf_ram.memory\[101\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__04845__A3 u_cpu.cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[30\]_D u_arbiter.i_wb_cpu_rdt\[27\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10195__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09233__A2 _04487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07244__A1 _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08441__B1 _04009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[45\] u_scanchain_local.module_data_in\[44\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[7\] u_scanchain_local.clk u_scanchain_local.module_data_in\[45\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__07795__A2 _03520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08992__A1 _04296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05528__B _01648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07547__A2 _03382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[16\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10119_ _00565_ io_in[4] u_cpu.rf_ram.memory\[136\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05653__S1 _01574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11099_ _11099_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_110_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05660_ _01542_ _02145_ _01418_ _02146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_90_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05591_ _02071_ _02073_ _02075_ _02077_ _01628_ _02078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__05730__A1 _02206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07330_ u_cpu.rf_ram.memory\[49\]\[3\] _03255_ _03259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10538__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06286__A2 _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07261_ _03220_ _00523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08680__B1 _04157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09000_ _04286_ _04359_ _04362_ _01121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06212_ _02475_ _02612_ _02613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09830__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07192_ _03169_ _03176_ _03182_ _00492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_u_scanchain_local.scan_flop\[21\]_D u_arbiter.i_wb_cpu_rdt\[18\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09224__A2 _04487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06038__A2 _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06143_ u_cpu.rf_ram.memory\[20\]\[2\] _02563_ _02566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10688__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07786__A2 _03520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06074_ _02522_ _02463_ _02523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05341__S0 _01646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05025_ _01445_ _01521_ _01522_ u_arbiter.o_wb_cpu_adr\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09902_ _00356_ io_in[4] u_cpu.rf_ram.memory\[60\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09980__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08735__A1 _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07538__A2 _03372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09833_ _00287_ io_in[4] u_cpu.rf_ram.memory\[67\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09764_ _00218_ io_in[4] u_cpu.rf_ram.memory\[119\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05644__S1 _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06976_ _02602_ _02684_ _03060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07145__S _03148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08468__C _03801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08715_ _04187_ _01011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_55_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05927_ _02375_ _02390_ _02407_ _02408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_09695_ _00149_ io_in[4] u_cpu.rf_ram.memory\[43\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10068__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09160__A1 _04284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05173__B _01654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05858_ u_cpu.cpu.genblk3.csr.mcause3_0\[0\] _02341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08646_ u_cpu.rf_ram.memory\[30\]\[4\] _04145_ _04150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07710__A2 _02638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05789_ u_cpu.rf_ram.memory\[92\]\[7\] u_cpu.rf_ram.memory\[93\]\[7\] u_cpu.rf_ram.memory\[94\]\[7\]
+ u_cpu.rf_ram.memory\[95\]\[7\] _01610_ _01611_ _02274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08577_ _04110_ _00950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07528_ _03371_ _03372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09463__A2 _04625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06277__A2 _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07459_ _03167_ _03325_ _03330_ _00611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10470_ _00903_ io_in[4] u_cpu.cpu.decode.op26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_u_scanchain_local.scan_flop\[12\]_D u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09215__A2 _04470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05580__S0 _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07226__A1 _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09129_ u_cpu.rf_ram.memory\[107\]\[4\] _04429_ _04434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07777__A2 _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[39\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05788__A1 _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05332__S0 _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07529__A2 _03372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11022_ _11022_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_104_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05635__S1 _01681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07055__S _03100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09703__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07701__A2 _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10806_ _01235_ io_in[4] u_cpu.rf_ram.memory\[85\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09853__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06268__A2 _02641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07465__A1 _03173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10737_ _01166_ io_in[4] u_cpu.rf_ram.memory\[105\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08662__B1 _04157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10830__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09206__A2 _04470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05102__I _01540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10668_ _01097_ io_in[4] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05571__S0 _01578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08265__I0 u_arbiter.i_wb_cpu_rdt\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07738__B _01369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10599_ _01028_ io_in[4] u_cpu.rf_ram.memory\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07768__A2 _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05323__S0 _01619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05258__B _01654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06440__A2 _02740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08568__I1 u_arbiter.i_wb_cpu_dbus_adr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09390__A1 _04191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05626__S1 _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06830_ _02967_ _02972_ _02979_ _00333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10210__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07940__A2 _03606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06761_ u_cpu.rf_ram.memory\[65\]\[3\] _02934_ _02938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05951__A1 _01403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09142__A1 _04284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05712_ u_cpu.rf_ram.memory\[68\]\[6\] u_cpu.rf_ram.memory\[69\]\[6\] u_cpu.rf_ram.memory\[70\]\[6\]
+ u_cpu.rf_ram.memory\[71\]\[6\] _01555_ _01652_ _02198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08500_ _03786_ _03860_ _03849_ _04061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09480_ _02590_ u_cpu.rf_ram.memory\[0\]\[4\] _04634_ _04639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06692_ _02899_ _00275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10360__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08431_ _03807_ _03809_ _04000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05643_ _01406_ _02080_ _02129_ _00005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_24_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08362_ _03876_ _03937_ _03938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05574_ u_cpu.rf_ram.memory\[52\]\[5\] u_cpu.rf_ram.memory\[53\]\[5\] u_cpu.rf_ram.memory\[54\]\[5\]
+ u_cpu.rf_ram.memory\[55\]\[5\] _01590_ _01591_ _02061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09445__A2 _04615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07313_ _03165_ _03245_ _03249_ _00546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06259__A2 _02641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08293_ u_cpu.rf_ram.memory\[114\]\[1\] _03879_ _03881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07244_ _03167_ _03206_ _03211_ _00515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05562__S0 _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07208__A1 _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07175_ _03171_ _03159_ _03172_ _00485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07759__A2 _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06126_ _02497_ _02551_ _02555_ _00053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05314__S0 _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06057_ _02477_ _02507_ _02508_ _00031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06431__A2 _02740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05008_ u_arbiter.i_wb_cpu_dbus_adr\[22\] _01442_ _01510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09726__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08479__B _03788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09381__A1 u_cpu.cpu.genblk3.csr.o_new_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09816_ _00270_ io_in[4] u_cpu.rf_ram.memory\[75\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05617__S1 _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07931__A2 _03596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[69\]_SI u_arbiter.o_wb_cpu_adr\[31\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_09747_ _00201_ io_in[4] u_cpu.rf_ram.memory\[17\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10703__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05942__A1 _02320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06959_ _03050_ _03051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09678_ _00132_ io_in[4] u_cpu.rf_ram.memory\[51\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09876__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07695__A1 _03343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08629_ _02372_ _02773_ _04138_ _04139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06498__A2 _02612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10853__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07447__A1 _03173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07998__A2 _03636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06018__I _02474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10522_ _00955_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10453_ _00886_ io_in[4] u_cpu.cpu.decode.opcode\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06670__A2 _02884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10384_ _00817_ io_in[4] u_cpu.rf_ram.memory\[122\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05305__S0 _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06422__A2 _02729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10233__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__04984__A2 _01442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11005_ _11005_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_42_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07922__A2 _03596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10383__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05933__A1 _02320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09124__A1 _04284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08609__S _04115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05541__B _01417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09427__A2 _04605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07989__A2 _03636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06110__A1 _02502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05290_ _01771_ _01780_ _01781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06661__A2 _02874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08402__A3 _03826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09749__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07610__A1 _03353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06413__A2 _02729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08980_ _04284_ _04349_ _04351_ _01112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07931_ u_cpu.rf_ram.memory\[112\]\[7\] _03596_ _03604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10726__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07862_ _03555_ _03558_ _03566_ _00779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09899__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09601_ _00055_ io_in[4] u_cpu.rf_ram.memory\[18\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08961__I1 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06813_ u_cpu.rf_ram.memory\[29\]\[7\] _02955_ _02970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05435__C _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07793_ u_cpu.rf_ram.memory\[34\]\[4\] _03520_ _03525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09532_ u_cpu.rf_ram.memory\[89\]\[3\] _04664_ _04668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06744_ _02746_ _02924_ _02928_ _00298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08519__S _01437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10876__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07677__A1 u_cpu.cpu.mem_bytecnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09463_ u_cpu.rf_ram.memory\[24\]\[4\] _04625_ _04630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06675_ u_cpu.rf_ram.memory\[75\]\[5\] _02884_ _02890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08414_ _03816_ _03979_ _03983_ _03984_ _00913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_05626_ u_cpu.rf_ram.memory\[72\]\[5\] u_cpu.rf_ram.memory\[73\]\[5\] u_cpu.rf_ram.memory\[74\]\[5\]
+ u_cpu.rf_ram.memory\[75\]\[5\] _01610_ _01611_ _02113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_40_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05152__A2 _01643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09394_ _04588_ _04589_ _04590_ _04591_ _01286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__05783__S0 _01619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10106__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07429__A1 _03173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05557_ _01542_ _02043_ _02044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08345_ _03921_ _03916_ _03922_ _03877_ _00906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_138_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08276_ _02343_ _03740_ _03866_ _00893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08254__S _01437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05488_ u_cpu.rf_ram.memory\[48\]\[4\] u_cpu.rf_ram.memory\[49\]\[4\] u_cpu.rf_ram.memory\[50\]\[4\]
+ u_cpu.rf_ram.memory\[51\]\[4\] _01544_ _01548_ _01976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_22_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05455__A3 _01943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06652__A2 _02874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07227_ u_cpu.rf_ram.memory\[70\]\[5\] _03196_ _03202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10256__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08929__A1 _04284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07158_ _02486_ _03161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06109_ u_cpu.rf_ram.memory\[81\]\[4\] _02541_ _02546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06404__A2 _02718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07089_ _02959_ _03119_ _03122_ _00449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05915__A1 _01374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09106__A1 _04284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07668__A1 _03357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05361__B _01565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05774__S0 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09409__A2 _04595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06891__A2 _03012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08391__C _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10505_ _00938_ io_in[4] u_cpu.rf_ram.memory\[31\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06643__A2 _02864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10436_ _00869_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10749__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08396__A2 u_arbiter.i_wb_cpu_rdt\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10367_ _00800_ io_in[4] u_cpu.rf_ram.memory\[11\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10298_ _00731_ io_in[4] u_cpu.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09345__A1 _04468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08148__A2 _03747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06159__A1 _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10899__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10129__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08320__A2 _03831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06460_ _02590_ u_cpu.rf_ram.memory\[4\]\[4\] _02756_ _02761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05765__S0 _01623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05411_ u_cpu.rf_ram.memory\[36\]\[3\] u_cpu.rf_ram.memory\[37\]\[3\] u_cpu.rf_ram.memory\[38\]\[3\]
+ u_cpu.rf_ram.memory\[39\]\[3\] _01619_ _01620_ _01900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_15_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06882__A2 _03002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06391_ _02482_ _02718_ _02719_ _00154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10279__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08130_ u_cpu.rf_ram.memory\[113\]\[3\] _03731_ _03735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05342_ _01645_ _01831_ _01648_ _01832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05517__S0 _01646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08061_ u_arbiter.i_wb_cpu_rdt\[10\] _03669_ _03678_ u_arbiter.i_wb_cpu_dbus_dat\[10\]
+ _03691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05273_ _01553_ _01763_ _01565_ _01764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06634__A2 _02864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07012_ _02524_ _02684_ _03080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08963_ u_arbiter.i_wb_cpu_rdt\[26\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[10\]
+ _04331_ _04342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__04948__A2 _01462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08139__A2 _03731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07914_ _03594_ _00803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08894_ _04290_ _04299_ _04304_ _01073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07845_ _02821_ _02893_ _03557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07898__A1 _02577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07776_ _03353_ _03510_ _03515_ _00744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04988_ _01445_ _01493_ _01494_ u_arbiter.o_wb_cpu_adr\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09515_ _04476_ _04654_ _04658_ _01340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08476__C _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06727_ u_cpu.rf_ram.memory\[67\]\[4\] _02914_ _02919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09446_ _04478_ _04615_ _04620_ _01309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06322__A1 _02502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06658_ _02750_ _02874_ _02880_ _00260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05756__S0 _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05609_ u_cpu.rf_ram.memory\[116\]\[5\] u_cpu.rf_ram.memory\[117\]\[5\] u_cpu.rf_ram.memory\[118\]\[5\]
+ u_cpu.rf_ram.memory\[119\]\[5\] _01623_ _01624_ _02096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_40_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09377_ _01381_ _01392_ _04568_ _04579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_40_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06873__A2 _03002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09914__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06589_ u_cpu.rf_ram.memory\[129\]\[7\] _02834_ _02842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04884__A1 _01408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08328_ _03773_ _03908_ _03909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08075__A1 u_arbiter.i_wb_cpu_rdt\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05508__S0 _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06625__A2 _02854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08259_ _03754_ _03800_ _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08378__A2 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10221_ _00667_ io_in[4] u_cpu.rf_ram.memory\[124\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10152_ _00598_ io_in[4] u_cpu.rf_ram.memory\[132\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09327__A1 _04468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05356__B _01654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10083_ _00529_ io_in[4] u_cpu.rf_ram.memory\[138\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06031__I _02486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08550__A2 _04094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06561__A1 _02744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07063__S _03100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10985_ _10985_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_16_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08302__A2 _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05091__B _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10421__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05747__S0 _01578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09594__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06864__A2 _02992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04875__A1 u_cpu.cpu.immdec.imm24_20\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10571__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06616__A2 _02854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05110__I _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10419_ _00852_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07041__A2 _03091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05960_ u_cpu.rf_ram_if.rdata0\[6\] _01403_ _02429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_04911_ _01433_ u_arbiter.o_wb_cpu_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05891_ _02361_ _02372_ _02373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_94_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08541__A2 _04084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07630_ _03355_ _03422_ _03428_ _00684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_04842_ u_cpu.cpu.bufreg.lsb\[0\] u_cpu.cpu.bufreg.lsb\[1\] u_arbiter.i_wb_cpu_dbus_sel\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_26_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06552__A1 _02754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07561_ u_cpu.rf_ram.memory\[126\]\[7\] _03382_ _03390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09937__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09300_ u_cpu.rf_ram.memory\[86\]\[5\] _04526_ _04532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06512_ u_cpu.rf_ram.memory\[16\]\[6\] _02791_ _02798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07492_ u_cpu.rf_ram.memory\[22\]\[2\] _03345_ _03350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[61\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05738__S0 _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09231_ u_cpu.rf_ram.memory\[59\]\[6\] _04487_ _04494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06855__A2 _02992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06443_ u_cpu.rf_ram.memory\[50\]\[5\] _02740_ _02751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10914__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09162_ _04286_ _04449_ _04452_ _01193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06374_ u_cpu.rf_ram.memory\[43\]\[1\] _02708_ _02710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07500__I _02506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05325_ u_cpu.rf_ram.memory\[32\]\[2\] u_cpu.rf_ram.memory\[33\]\[2\] u_cpu.rf_ram.memory\[34\]\[2\]
+ u_cpu.rf_ram.memory\[35\]\[2\] _01623_ _01624_ _01815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08113_ _03723_ _03718_ _03724_ _00872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07804__A1 _03343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06607__A2 _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09093_ u_cpu.rf_ram.memory\[105\]\[4\] _04409_ _04414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05256_ _01541_ _01746_ _01747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08044_ _03677_ _03679_ _00848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07280__A2 _03225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05291__A1 _01406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09557__A1 _04482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05830__A3 _02313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05187_ _01657_ _01678_ _01402_ _01679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07032__A2 _03091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09995_ _00002_ io_in[4] u_cpu.rf_ram.rdata\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09309__A1 _04468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08946_ _04333_ _01096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05433__I3 u_cpu.rf_ram.memory\[119\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[14\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06918__I0 _02596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08877_ _02511_ _04294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08532__A2 _04084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10444__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07828_ u_cpu.rf_ram.memory\[120\]\[2\] _03541_ _03546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05346__A2 _01835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07759_ u_cpu.rf_ram.memory\[92\]\[5\] _03500_ _03506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08296__A1 _03545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07099__A2 _03119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[29\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10770_ _01199_ io_in[4] u_cpu.rf_ram.memory\[69\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10594__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09429_ u_cpu.rf_ram.memory\[26\]\[5\] _04605_ _04611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06846__A2 _02982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04857__A1 _01369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08048__A1 u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08048__B2 u_arbiter.i_wb_cpu_dbus_dat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05806__B1 _02288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07271__A2 _03225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05282__A1 _01399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10204_ _00650_ io_in[4] u_cpu.rf_ram.memory\[126\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07023__A2 _03081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10135_ _00581_ io_in[4] u_cpu.rf_ram.memory\[134\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06782__A1 _02748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10066_ _00512_ io_in[4] u_cpu.rf_ram.memory\[143\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08523__A2 _02448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05533__C _01426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10937__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08287__A1 _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10968_ _10968_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__08287__B2 _03876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08617__S _04115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05105__I _01397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06837__A2 _02982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10899_ _01328_ io_in[4] u_cpu.rf_ram.memory\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08039__A1 _02781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05110_ _01543_ _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06090_ u_cpu.rf_ram.memory\[21\]\[4\] _02530_ _02535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10317__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05273__A1 _01553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09539__A1 _04482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05041_ _01443_ _01533_ _01534_ u_arbiter.o_wb_cpu_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08211__A1 _03776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07014__A2 _03081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05025__A1 _01445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08800_ _02433_ _02453_ _04236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_140_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10467__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09780_ _00234_ io_in[4] u_cpu.rf_ram.memory\[139\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06992_ u_cpu.rf_ram.memory\[55\]\[7\] _03061_ _03069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05120__S1 _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08731_ _04198_ _04199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05943_ _02320_ _02418_ _02419_ _00018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_26_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08662_ u_cpu.cpu.ctrl.o_ibus_adr\[2\] _04155_ _04157_ u_cpu.cpu.ctrl.o_ibus_adr\[3\]
+ _04160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__05724__B _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05874_ u_cpu.cpu.state.o_cnt_r\[0\] _02338_ _02356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06525__A1 _02746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07613_ u_cpu.rf_ram.memory\[123\]\[6\] _03412_ _03419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08593_ u_arbiter.i_wb_cpu_dbus_adr\[17\] u_arbiter.i_wb_cpu_dbus_adr\[16\] _04115_
+ _04119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_35_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07544_ _03359_ _03372_ _03380_ _00646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08278__A1 _03801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06828__A2 _02972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07475_ _02590_ u_cpu.rf_ram.memory\[12\]\[4\] _03334_ _03339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09214_ _02516_ _04484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06426_ _02469_ _02684_ _02739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09145_ u_cpu.rf_ram.memory\[83\]\[3\] _04439_ _04443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06357_ u_cpu.rf_ram.memory\[41\]\[2\] _02697_ _02700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05308_ _01542_ _01797_ _01418_ _01798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06288_ _02512_ _02651_ _02658_ _00112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09076_ _04290_ _04399_ _04404_ _01155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08450__B2 _03855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05264__A1 _01645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08027_ u_arbiter.i_wb_cpu_dbus_dat\[2\] _03658_ _03665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05239_ _01723_ _01725_ _01727_ _01729_ _01628_ _01730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_116_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07005__A2 _03071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08202__A1 _03773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09250__I0 _02599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09978_ _00432_ io_in[4] u_cpu.rf_ram.memory\[9\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06764__A1 _02748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08929_ _04284_ _04322_ _04324_ _01088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08505__A2 _04016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06516__A1 _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10822_ _01251_ io_in[4] u_cpu.rf_ram.memory\[86\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08269__A1 _03767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10753_ _01182_ io_in[4] u_cpu.rf_ram.memory\[107\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06819__A2 _02972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10684_ _01113_ io_in[4] u_cpu.rf_ram.memory\[101\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07492__A2 _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09632__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08441__A1 _03744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08172__S _01435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07244__A2 _03206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08441__B2 _03876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08992__A2 _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[38\] u_scanchain_local.module_data_in\[37\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[0\] u_scanchain_local.clk u_scanchain_local.module_data_in\[38\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_5_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09782__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08744__A2 _04199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10118_ _00564_ io_in[4] u_cpu.rf_ram.memory\[136\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11098_ _11098_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05544__B _01402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__04939__I _01442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10049_ _00495_ io_in[4] u_cpu.rf_ram.memory\[71\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06507__A1 _02746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05590_ _01645_ _02076_ _01626_ _02077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05730__A2 _02215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07260_ _02590_ u_cpu.rf_ram.memory\[14\]\[4\] _03215_ _03220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06211_ _02464_ _02560_ _02612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07191_ u_cpu.rf_ram.memory\[73\]\[5\] _03176_ _03182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06142_ _02487_ _02563_ _02565_ _00059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09480__I0 _02590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07235__A2 _03206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08983__A2 _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06073_ _02456_ _02458_ _02522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__05341__S1 _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05797__A2 _02277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06994__A1 _02684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05024_ u_arbiter.i_wb_cpu_dbus_adr\[26\] _01457_ _01522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09901_ _00355_ io_in[4] u_cpu.rf_ram.memory\[60\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08735__A2 _04199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09832_ _00286_ io_in[4] u_cpu.rf_ram.memory\[68\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06746__A1 _02748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09763_ _00217_ io_in[4] u_cpu.rf_ram.memory\[119\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06975_ _02969_ _03051_ _03059_ _00398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08714_ u_cpu.cpu.ctrl.o_ibus_adr\[27\] _04173_ _04175_ u_cpu.cpu.ctrl.o_ibus_adr\[28\]
+ _04187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08499__A1 _03742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04849__I _01374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05926_ _01374_ _02391_ _02406_ _02407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_39_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09694_ _00148_ io_in[4] u_cpu.rf_ram.memory\[43\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09160__A2 _04449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08645_ _03547_ _04145_ _04149_ _00979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05857_ _02337_ u_cpu.cpu.state.o_cnt_r\[3\] _02338_ _02339_ _02340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_15_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08576_ u_arbiter.i_wb_cpu_dbus_adr\[9\] u_arbiter.i_wb_cpu_dbus_adr\[8\] _02445_
+ _04110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05788_ _01422_ _02263_ _02272_ _02273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_74_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08484__C _03797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07527_ _02727_ _02821_ _03371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08120__B1 _03718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09655__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07458_ u_cpu.rf_ram.memory\[130\]\[4\] _03325_ _03330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06409_ u_cpu.rf_ram.memory\[47\]\[0\] _02729_ _02730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07389_ _03169_ _03285_ _03291_ _00580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05580__S1 _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09128_ _04288_ _04429_ _04433_ _01178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10632__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07226__A2 _03196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09059_ u_cpu.rf_ram.memory\[99\]\[5\] _04389_ _04395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05629__B _01417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05332__S1 _01616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05788__A2 _02263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06985__A1 _02961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08005__B u_cpu.cpu.mem_bytecnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10782__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11021_ _11021_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_104_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[7\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10012__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05960__A2 _01403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09151__A2 _04439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10162__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10805_ _01234_ io_in[4] u_cpu.rf_ram.memory\[85\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10736_ _01165_ io_in[4] u_cpu.rf_ram.memory\[105\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07465__A2 _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10667_ _01096_ io_in[4] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05571__S1 _01580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08414__A1 _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07217__A2 _03196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08265__I1 u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10598_ _01027_ io_in[4] u_cpu.rf_ram.memory\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07738__C _01370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06976__A1 _02602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05323__S1 _01620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06728__A1 _02748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09390__A2 _02348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06760_ _02744_ _02934_ _02937_ _00305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09142__A2 _04439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05711_ _01667_ _02196_ _02197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10505__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06691_ _02590_ u_cpu.rf_ram.memory\[6\]\[4\] _02894_ _02899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08430_ _02765_ u_arbiter.i_wb_cpu_rdt\[7\] _03998_ _03999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05642_ _02119_ _02128_ _02129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09678__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06900__A1 _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08361_ _03755_ _03757_ _03780_ _03936_ _03937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05573_ _02053_ _02055_ _02057_ _02059_ _01426_ _02060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_108_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07312_ u_cpu.rf_ram.memory\[137\]\[3\] _03245_ _03249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10655__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08292_ _03539_ _03879_ _03880_ _00895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07456__A2 _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08653__A1 _03555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05467__A1 _01406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07243_ u_cpu.rf_ram.memory\[143\]\[4\] _03206_ _03211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05562__S1 _01557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07208__A2 _03186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07174_ u_cpu.rf_ram.memory\[72\]\[6\] _03159_ _03172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06125_ u_cpu.rf_ram.memory\[18\]\[3\] _02551_ _02555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05449__B _01565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05609__I3 u_cpu.rf_ram.memory\[119\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05314__S1 _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06967__A1 _02961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06056_ u_cpu.rf_ram.memory\[82\]\[5\] _02477_ _02508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05007_ _01506_ _01507_ _01509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08708__A2 _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10035__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09815_ _00269_ io_in[4] u_cpu.rf_ram.memory\[75\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09746_ _00200_ io_in[4] u_cpu.rf_ram.memory\[17\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05184__B _01417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06958_ _02684_ _02810_ _03050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09371__S _04568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09133__A2 _04429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10185__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05909_ _02381_ _02382_ _02347_ _02389_ _02390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_55_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09677_ _00131_ io_in[4] u_cpu.rf_ram.memory\[51\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06889_ u_cpu.rf_ram.memory\[19\]\[0\] _03012_ _03013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08628_ u_cpu.cpu.state.o_cnt_r\[0\] u_cpu.cpu.state.o_cnt_r\[1\] _02338_ _02773_
+ _04138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__06794__I _02486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07695__A2 _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08892__A1 _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[0\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08559_ _03553_ _04094_ _04101_ _00941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07447__A2 _03315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05458__A1 _01399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10521_ _00954_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10452_ _00885_ io_in[4] u_cpu.cpu.decode.opcode\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10383_ _00816_ io_in[4] u_cpu.rf_ram.memory\[122\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06958__A1 _02684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05305__S1 _01574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05481__I1 u_cpu.rf_ram.memory\[29\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07066__S _03109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11004_ _11004_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_120_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08389__C _03800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10528__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05806__C _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07383__A1 _03163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09820__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09124__A2 _04429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07135__A1 _02969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10678__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08883__A1 _02475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09970__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08635__A1 _02431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07438__A2 _03315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05113__I _01416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05449__A1 _01553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10719_ _01148_ io_in[4] u_cpu.rf_ram.memory\[99\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06110__A2 _02541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08938__A2 _04322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09060__A1 _04292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10058__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06949__A1 _02961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07610__A2 _03412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07930_ _03553_ _03596_ _03603_ _00810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07861_ u_cpu.rf_ram.memory\[118\]\[7\] _03558_ _03566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09600_ _00054_ io_in[4] u_cpu.rf_ram.memory\[18\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06812_ _02516_ _02969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07792_ _03351_ _03520_ _03524_ _00751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09531_ _04474_ _04664_ _04667_ _01347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09115__A2 _04419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06743_ u_cpu.rf_ram.memory\[66\]\[3\] _02924_ _02928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09462_ _04476_ _04625_ _04629_ _01316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06674_ _02748_ _02884_ _02889_ _00267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_u_scanchain_local.scan_flop\[29\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07677__A2 _03454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07503__I _02511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08413_ u_cpu.cpu.immdec.imm30_25\[4\] _03949_ _03976_ u_cpu.cpu.immdec.imm30_25\[5\]
+ _03984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_05625_ _01553_ _02111_ _01565_ _02112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09393_ u_cpu.cpu.genblk3.csr.mstatus_mie _04565_ _04590_ _04591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_40_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05783__S1 _01620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08344_ u_cpu.cpu.immdec.imm24_20\[3\] _03914_ _03797_ _03922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05556_ u_cpu.rf_ram.memory\[8\]\[5\] u_cpu.rf_ram.memory\[9\]\[5\] u_cpu.rf_ram.memory\[10\]\[5\]
+ u_cpu.rf_ram.memory\[11\]\[5\] _01546_ _01550_ _02043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_33_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07429__A2 _03305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08275_ _03816_ _03856_ _03865_ _02768_ _03866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06101__A2 _02541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05487_ _01589_ _01974_ _01975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07226_ _03167_ _03196_ _03201_ _00507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08929__A2 _04322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07157_ _03157_ _03159_ _03160_ _00479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06108_ _02497_ _02541_ _02545_ _00045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07601__A2 _03412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07088_ u_cpu.rf_ram.memory\[142\]\[2\] _03119_ _03122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05612__A1 _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06039_ _02477_ _02492_ _02493_ _00028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06789__I _02481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09843__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09354__A2 _04556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07365__A1 _03163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10820__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05915__A2 _02391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09106__A2 _04419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09729_ _00183_ io_in[4] u_cpu.rf_ram.memory\[4\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07117__A1 _02969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09993__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07668__A2 _03442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06340__A2 _02686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05774__S1 _01549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08093__A2 _03683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10200__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10504_ _00937_ io_in[4] u_cpu.rf_ram.memory\[31\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07840__A2 _03541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05851__A1 _02332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10435_ _00868_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09042__A1 _04292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10366_ _00799_ io_in[4] u_cpu.rf_ram.memory\[11\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10350__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xu_scanchain_local.scan_flop\[20\] u_arbiter.i_wb_cpu_rdt\[17\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[14\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10297_ _00730_ io_in[4] u_cpu.cpu.bufreg2.i_cnt_done vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09345__A2 _04556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06159__A2 _01386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08156__I0 u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05552__B _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08856__A1 _03555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07659__A2 _03442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07903__I0 _02584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05765__S1 _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05410_ _01614_ _01898_ _01605_ _01899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06390_ u_cpu.rf_ram.memory\[48\]\[0\] _02718_ _02719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05341_ u_cpu.rf_ram.memory\[120\]\[2\] u_cpu.rf_ram.memory\[121\]\[2\] u_cpu.rf_ram.memory\[122\]\[2\]
+ u_cpu.rf_ram.memory\[123\]\[2\] _01646_ _01603_ _01831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__04893__A2 _01368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09281__A1 _04478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09716__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05517__S1 _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06095__A1 _02512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08060_ u_arbiter.i_wb_cpu_dbus_dat\[11\] _03683_ _03690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05272_ u_cpu.rf_ram.memory\[68\]\[1\] u_cpu.rf_ram.memory\[69\]\[1\] u_cpu.rf_ram.memory\[70\]\[1\]
+ u_cpu.rf_ram.memory\[71\]\[1\] _01555_ _01652_ _01763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07831__A2 _03541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07011_ _02969_ _03071_ _03079_ _00414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09866__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06398__A2 _02718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08962_ _04341_ _01104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10843__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09336__A2 _04546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07913_ _02599_ u_cpu.rf_ram.memory\[11\]\[7\] _03586_ _03594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_64_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08893_ u_cpu.rf_ram.memory\[95\]\[4\] _04299_ _04304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07347__A1 _03163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07844_ _03555_ _03541_ _03556_ _00771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07898__A2 _02706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07775_ u_cpu.rf_ram.memory\[35\]\[4\] _03510_ _03515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04987_ u_arbiter.i_wb_cpu_dbus_adr\[17\] _01457_ _01494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06570__A2 _02823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09514_ u_cpu.rf_ram.memory\[100\]\[3\] _04654_ _04658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06726_ _02746_ _02914_ _02918_ _00290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09445_ u_cpu.rf_ram.memory\[25\]\[4\] _04615_ _04620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06657_ u_cpu.rf_ram.memory\[76\]\[5\] _02874_ _02880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06322__A2 _02673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10223__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05756__S1 _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05608_ _01541_ _02094_ _02095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08265__S _01437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09376_ u_cpu.cpu.genblk3.csr.mcause3_0\[3\] _04578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06588_ _02752_ _02834_ _02841_ _00229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04884__A2 _01409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08327_ _03763_ _03860_ _03828_ _03744_ _03800_ _03908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_138_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05539_ _01667_ _02026_ _02027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08075__A2 _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05508__S1 _01616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08258_ _03773_ _03848_ _03849_ _03850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__07822__A2 _03541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10373__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05833__A1 _01369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07209_ u_cpu.rf_ram.memory\[71\]\[5\] _03186_ _03192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09024__A1 _04292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08189_ _03745_ _03788_ _03789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_10220_ _00666_ io_in[4] u_cpu.rf_ram.memory\[124\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07586__A1 _03347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10151_ _00597_ io_in[4] u_cpu.rf_ram.memory\[132\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09327__A2 _04546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10082_ _00528_ io_in[4] u_cpu.rf_ram.memory\[138\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06561__A2 _02823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05372__B _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10984_ _10984_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_43_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09739__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06313__A2 _02673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05747__S1 _01580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08175__S _01435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04875__A2 _01388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10716__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09263__A1 _04478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08066__A2 _03683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[68\] u_scanchain_local.module_data_in\[67\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[30\] u_scanchain_local.clk u_scanchain_local.module_data_in\[68\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_11_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09889__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07813__A2 _03530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05824__A1 _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10866__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10418_ _00851_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10349_ _00782_ io_in[4] u_cpu.rf_ram.memory\[121\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09318__A2 _04536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07329__A1 _03163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04910_ u_arbiter.i_wb_cpu_ibus_adr\[1\] _01431_ _01433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_39_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05890_ _02371_ _02372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07254__S _03215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06001__A1 _02312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04841_ _01368_ u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06552__A2 _02812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10246__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07560_ _03357_ _03382_ _03389_ _00653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08829__A1 u_cpu.cpu.immdec.imm11_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06511_ _02750_ _02791_ _02797_ _00196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07491_ _02491_ _03349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06304__A2 _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07501__A1 u_cpu.rf_ram.memory\[22\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05738__S1 _01557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09230_ _04480_ _04487_ _04493_ _01220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06442_ _02506_ _02750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10396__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09161_ u_cpu.rf_ram.memory\[108\]\[2\] _04449_ _04452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06373_ _02482_ _02708_ _02709_ _00146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08057__A2 _03683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08112_ u_arbiter.i_wb_cpu_rdt\[28\] _03653_ _03654_ u_arbiter.i_wb_cpu_dbus_dat\[28\]
+ _03724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05324_ _01589_ _01813_ _01814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09092_ _04288_ _04409_ _04413_ _01162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07804__A2 _03530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08043_ u_arbiter.i_wb_cpu_rdt\[4\] _03669_ _03678_ u_arbiter.i_wb_cpu_dbus_dat\[4\]
+ _03679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05255_ u_cpu.rf_ram.memory\[112\]\[1\] u_cpu.rf_ram.memory\[113\]\[1\] u_cpu.rf_ram.memory\[114\]\[1\]
+ u_cpu.rf_ram.memory\[115\]\[1\] _01590_ _01591_ _01746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09006__A1 _04292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05291__A2 _01732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09557__A2 _04674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05186_ _01539_ _01666_ _01677_ _01678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__07568__A1 _03347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09994_ _00001_ io_in[4] u_cpu.rf_ram.rdata\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09309__A2 _04536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08945_ u_arbiter.i_wb_cpu_rdt\[17\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\]
+ _04331_ _04333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_9_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08876_ _04292_ _04282_ _04293_ _01066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07827_ _02491_ _03545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06543__A2 _02812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07740__A1 _02333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07758_ _03353_ _03500_ _03505_ _00736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_77_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06709_ u_cpu.rf_ram.memory\[68\]\[4\] _02904_ _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10739__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09493__A1 _04472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08296__A2 _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07689_ _01428_ _02376_ _00709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_44_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09428_ _04478_ _04605_ _04610_ _01301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04857__A2 _01370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09359_ _04484_ _04556_ _04564_ _01278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08048__A2 _03653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06059__A1 _02460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10889__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05657__I1 u_cpu.rf_ram.memory\[29\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05282__A2 _01772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09548__A2 _04674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10119__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10203_ _00649_ io_in[4] u_cpu.rf_ram.memory\[126\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10134_ _00580_ io_in[4] u_cpu.rf_ram.memory\[134\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08359__I0 u_arbiter.i_wb_cpu_rdt\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06782__A2 _02944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10269__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10065_ _00511_ io_in[4] u_cpu.rf_ram.memory\[143\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07074__S _03109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10967_ _10967_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_91_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08287__A2 _03867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10898_ _01327_ io_in[4] u_cpu.rf_ram.memory\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08039__A2 _03648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07798__A1 _03357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09539__A2 _04664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06470__A1 _02765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05040_ u_arbiter.i_wb_cpu_dbus_adr\[30\] _01457_ _01534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05277__B _01417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08211__A2 _03768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06991_ _02967_ _03061_ _03068_ _00405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06773__A2 _02944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08730_ _02660_ _04197_ _04198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09904__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05942_ _02320_ u_cpu.rf_ram_if.rdata1\[4\] _02419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08661_ _04159_ _00985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_22_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05873_ u_cpu.cpu.alu.cmp_r _02355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_26_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05328__A3 _01817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06525__A2 _02801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07612_ _03355_ _03412_ _03418_ _00676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08770__I0 _02584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08592_ _04118_ _00957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07543_ u_cpu.rf_ram.memory\[127\]\[7\] _03372_ _03380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07474_ _03338_ _00618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09213_ _04482_ _04470_ _04483_ _01213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06425_ _02481_ _02738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09144_ _04286_ _04439_ _04442_ _01185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06356_ _02487_ _02697_ _02699_ _00139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05307_ u_cpu.rf_ram.memory\[24\]\[2\] u_cpu.rf_ram.memory\[25\]\[2\] u_cpu.rf_ram.memory\[26\]\[2\]
+ u_cpu.rf_ram.memory\[27\]\[2\] _01578_ _01580_ _01797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09075_ u_cpu.rf_ram.memory\[79\]\[4\] _04399_ _04404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06287_ u_cpu.rf_ram.memory\[46\]\[6\] _02651_ _02658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08450__A2 _04016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05264__A2 _01754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08026_ _03648_ _03663_ _03664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05238_ _01541_ _01728_ _01626_ _01729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_122_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05187__B _01402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05169_ _01645_ _01660_ _01648_ _01661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08202__A2 _03800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10411__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05016__A2 _01457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09977_ _00431_ io_in[4] u_cpu.rf_ram.memory\[9\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09584__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06764__A2 _02934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06797__I _02491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08928_ u_cpu.rf_ram.memory\[28\]\[1\] _04322_ _04324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08859_ _04281_ _04282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10561__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07713__A1 _03343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06516__A2 _02539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08761__I0 _02596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10821_ _01250_ io_in[4] u_cpu.rf_ram.memory\[86\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09466__A1 _04480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08269__A2 _03768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10752_ _01181_ io_in[4] u_cpu.rf_ram.memory\[107\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10683_ _01112_ io_in[4] u_cpu.rf_ram.memory\[101\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06037__I _02491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08441__A2 _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09927__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10091__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07252__I0 _02573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[60\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10904__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06755__A2 _02934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10117_ _00563_ io_in[4] u_cpu.rf_ram.memory\[136\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11097_ _11097_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_110_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10048_ _00494_ io_in[4] u_cpu.rf_ram.memory\[73\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06507__A2 _02791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05191__A1 _01399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[62\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08680__A2 _04155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06210_ _02611_ _00081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07190_ _03167_ _03176_ _03181_ _00491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06141_ u_cpu.rf_ram.memory\[20\]\[1\] _02563_ _02565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_u_scanchain_local.scan_flop\[13\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08432__A2 _03831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10434__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06072_ _02467_ _02520_ _02521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_104_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06994__A2 _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05023_ u_cpu.cpu.ctrl.o_ibus_adr\[26\] _01520_ _01521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09900_ _00354_ io_in[4] u_cpu.rf_ram.memory\[60\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08196__A1 _02765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[28\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09831_ _00285_ io_in[4] u_cpu.rf_ram.memory\[68\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10584__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06746__A2 _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05735__B _01417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09762_ _00216_ io_in[4] u_cpu.rf_ram.memory\[119\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06974_ u_cpu.rf_ram.memory\[56\]\[7\] _03051_ _03059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07506__I _02516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05925_ _02404_ _02356_ _02405_ _02406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_39_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08713_ _04186_ _01010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_132_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09693_ _00147_ io_in[4] u_cpu.rf_ram.memory\[43\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05454__C _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08644_ u_cpu.rf_ram.memory\[30\]\[3\] _04145_ _04149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05856_ u_cpu.cpu.decode.op26 _01411_ _02339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_54_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07171__A2 _03159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08575_ _04109_ _00949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05182__A1 _01667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05787_ _02265_ _02267_ _02269_ _02271_ _01607_ _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__09448__A1 _04480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07526_ _03359_ _03362_ _03370_ _00638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08120__A1 u_arbiter.i_wb_cpu_rdt\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08120__B2 _02325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07457_ _03165_ _03325_ _03329_ _00610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06408_ _02728_ _02729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06682__A1 _02577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07388_ u_cpu.rf_ram.memory\[134\]\[5\] _03285_ _03291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09127_ u_cpu.rf_ram.memory\[107\]\[3\] _04429_ _04433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06339_ _02492_ _02686_ _02689_ _00132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09058_ _04290_ _04389_ _04394_ _01147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05788__A3 _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08005__C u_cpu.cpu.bufreg.lsb\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08009_ u_arbiter.i_wb_cpu_dbus_dat\[0\] _02774_ _03649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06985__A2 _03061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10927__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04996__A1 _01443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08187__A1 _03776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11020_ _11020_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_103_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06737__A2 _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08021__B _02781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07162__A2 _03159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10307__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05173__A1 _01553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10804_ _01233_ io_in[4] u_cpu.rf_ram.memory\[85\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10735_ _01164_ io_in[4] u_cpu.rf_ram.memory\[105\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08662__A2 _04155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10457__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10666_ _01095_ io_in[4] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_scanchain_local.scan_flop\[50\] u_scanchain_local.module_data_in\[49\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[12\] u_scanchain_local.clk u_scanchain_local.module_data_in\[50\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
X_10597_ _01026_ io_in[4] u_cpu.rf_ram.memory\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07473__I0 _02587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06976__A2 _02684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08178__A1 _02765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06728__A2 _02914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08973__I0 u_arbiter.i_wb_cpu_rdt\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05710_ u_cpu.rf_ram.memory\[64\]\[6\] u_cpu.rf_ram.memory\[65\]\[6\] u_cpu.rf_ram.memory\[66\]\[6\]
+ u_cpu.rf_ram.memory\[67\]\[6\] _01571_ _01668_ _02196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_110_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06690_ _02898_ _00274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07262__S _03215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08350__A1 _03742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05641_ _02121_ _02123_ _02125_ _02127_ _01404_ _02128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__05164__B2 _01655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06900__A2 _03012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08360_ _03741_ _03778_ _03779_ _03935_ _03936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08157__I _03756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05572_ _01542_ _02058_ _01418_ _02059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_32_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07311_ _03163_ _03245_ _03248_ _00545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08291_ u_cpu.rf_ram.memory\[114\]\[0\] _03879_ _03880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08653__A2 _04145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07242_ _03165_ _03206_ _03210_ _00514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05467__A2 _01906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07173_ _02511_ _03171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06416__A1 _02497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06124_ _02492_ _02551_ _02554_ _00052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06967__A2 _03051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06055_ _02506_ _02507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__04978__A1 u_cpu.cpu.ctrl.o_ibus_adr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08169__A1 _03767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05006_ _01506_ _01507_ _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_120_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06719__A2 _02914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09814_ _00268_ io_in[4] u_cpu.rf_ram.memory\[75\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07392__A2 _03285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09745_ _00199_ io_in[4] u_cpu.rf_ram.memory\[17\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06957_ _02969_ _03041_ _03049_ _00390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05908_ _01373_ _02383_ _00728_ _02388_ _02389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_28_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06888_ _03011_ _03012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09676_ _00130_ io_in[4] u_cpu.rf_ram.memory\[51\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09622__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08341__A1 u_cpu.cpu.immdec.imm24_20\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08627_ _04133_ _04135_ _04137_ _02445_ _00973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_05839_ u_cpu.rf_ram_if.rdata1\[0\] _02320_ _02323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08892__A2 _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__04902__A1 _01399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08558_ u_cpu.rf_ram.memory\[31\]\[6\] _04094_ _04101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07509_ _02612_ _02832_ _03361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08489_ _03743_ _03776_ _03779_ _04050_ _03851_ _04051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__09772__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08644__A2 _04145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10520_ _00953_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05458__A2 _01946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10451_ _00884_ io_in[4] u_cpu.cpu.decode.opcode\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06407__A1 _02639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10382_ _00815_ io_in[4] u_cpu.rf_ram.memory\[122\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06958__A2 _02810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05630__A2 _02112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11003_ _11003_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__08955__I0 u_arbiter.i_wb_cpu_rdt\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07383__A2 _03285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05394__A1 _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07135__A2 _03139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05146__A1 _01636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08883__A2 _02727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06894__A1 _02959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10718_ _01147_ io_in[4] u_cpu.rf_ram.memory\[99\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10649_ _01078_ io_in[4] u_cpu.rf_ram.memory\[96\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05269__C _01426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09060__A2 _04389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06949__A2 _03041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07860_ _03553_ _03558_ _03565_ _00778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09645__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09472__S _04634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07374__A2 _03275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06811_ _02967_ _02955_ _02968_ _00325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07791_ u_cpu.rf_ram.memory\[34\]\[3\] _03520_ _03524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05385__A1 _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09530_ u_cpu.rf_ram.memory\[89\]\[2\] _04664_ _04667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06742_ _02744_ _02924_ _02927_ _00297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10622__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08323__A1 _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07126__A2 _03139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09461_ u_cpu.rf_ram.memory\[24\]\[3\] _04625_ _04629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06673_ u_cpu.rf_ram.memory\[75\]\[4\] _02884_ _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05137__B2 _01627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09795__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08412_ _03927_ _03980_ _03982_ _03853_ _03983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_05624_ u_cpu.rf_ram.memory\[68\]\[5\] u_cpu.rf_ram.memory\[69\]\[5\] u_cpu.rf_ram.memory\[70\]\[5\]
+ u_cpu.rf_ram.memory\[71\]\[5\] _01555_ _01652_ _02111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09392_ _04191_ _02340_ _04590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08343_ u_cpu.cpu.immdec.imm24_20\[2\] _03921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_71_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05555_ _01406_ _01993_ _02042_ _00004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10772__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08626__A2 _02773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[6\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08274_ _03780_ _03857_ _03864_ _03865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05486_ u_cpu.rf_ram.memory\[52\]\[4\] u_cpu.rf_ram.memory\[53\]\[4\] u_cpu.rf_ram.memory\[54\]\[4\]
+ u_cpu.rf_ram.memory\[55\]\[4\] _01590_ _01591_ _01974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_20_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07225_ u_cpu.rf_ram.memory\[70\]\[4\] _03196_ _03201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10002__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07156_ u_cpu.rf_ram.memory\[72\]\[0\] _03159_ _03160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09051__A2 _04389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06107_ u_cpu.rf_ram.memory\[81\]\[3\] _02541_ _02545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07087_ _02957_ _03119_ _03121_ _00448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05612__A2 _02089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06038_ u_cpu.rf_ram.memory\[82\]\[2\] _02477_ _02493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10152__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07365__A2 _03275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05376__A1 _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07989_ u_cpu.rf_ram.memory\[33\]\[0\] _03636_ _03637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09728_ _00182_ io_in[4] u_cpu.rf_ram.memory\[4\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08314__A1 _03890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07117__A2 _03129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09659_ _00113_ io_in[4] u_cpu.rf_ram.memory\[46\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06876__A1 _02959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08078__B1 _03678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09290__A2 _04526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10503_ _00936_ io_in[4] u_cpu.rf_ram.memory\[31\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10434_ _00867_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05851__A2 _02333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09042__A2 _04379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08250__B1 _03818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10365_ _00798_ io_in[4] u_cpu.rf_ram.memory\[11\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09668__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10296_ _00729_ io_in[4] u_cpu.cpu.ctrl.i_jump vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05817__C _01404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_scanchain_local.scan_flop\[13\] u_arbiter.i_wb_cpu_rdt\[10\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[7\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_120_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10645__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07356__A2 _03265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08553__A1 _03547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05367__A1 _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07108__A2 _03129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10795__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08856__A2 _04271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05124__I _01547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10025__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05340_ _01398_ _01829_ _01830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09281__A2 _04516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05271_ _01667_ _01761_ _01762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07292__A1 u_cpu.rf_ram.memory\[39\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06095__A2 _02530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07010_ u_cpu.rf_ram.memory\[54\]\[7\] _03071_ _03079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05842__A2 _02325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10175__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09033__A2 _04379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07595__A2 _03402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08961_ u_arbiter.i_wb_cpu_rdt\[25\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[9\]
+ _04331_ _04341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07912_ _03593_ _00802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08892_ _04288_ _04299_ _04303_ _01072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07347__A2 _03265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08544__A1 _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07843_ u_cpu.rf_ram.memory\[120\]\[7\] _03541_ _03556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07774_ _03351_ _03510_ _03514_ _00743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_04986_ u_cpu.cpu.ctrl.o_ibus_adr\[17\] _01491_ _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_84_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09513_ _04474_ _04654_ _04657_ _01339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06725_ u_cpu.rf_ram.memory\[67\]\[3\] _02914_ _02918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08847__A2 _04271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06858__A1 _02959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06656_ _02748_ _02874_ _02879_ _00259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09444_ _04476_ _04615_ _04619_ _01308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05607_ u_cpu.rf_ram.memory\[112\]\[5\] u_cpu.rf_ram.memory\[113\]\[5\] u_cpu.rf_ram.memory\[114\]\[5\]
+ u_cpu.rf_ram.memory\[115\]\[5\] _01619_ _01620_ _02094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05530__A1 _01609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09375_ _04568_ _04576_ _04577_ _01281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06587_ u_cpu.rf_ram.memory\[129\]\[6\] _02834_ _02841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05538_ u_cpu.rf_ram.memory\[72\]\[4\] u_cpu.rf_ram.memory\[73\]\[4\] u_cpu.rf_ram.memory\[74\]\[4\]
+ u_cpu.rf_ram.memory\[75\]\[4\] _01610_ _01611_ _02026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08326_ _03895_ _03905_ _03906_ _03907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__04873__I _01398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09272__A2 _04516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10518__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08257_ _03786_ _03790_ _03831_ _03849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07283__A1 _03171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06086__A2 _02530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05469_ _01542_ _01956_ _01957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07208_ _03167_ _03186_ _03191_ _00499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05833__A2 _01372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08188_ u_arbiter.i_wb_cpu_rdt\[8\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[8\]
+ _01435_ _03788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09810__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09024__A2 _04369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07035__A1 _02957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07139_ _02581_ u_cpu.rf_ram.memory\[13\]\[1\] _03148_ _03150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_133_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10668__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07586__A2 _03402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10150_ _00596_ io_in[4] u_cpu.rf_ram.memory\[132\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05597__A1 _01594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09960__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10081_ _00527_ io_in[4] u_cpu.rf_ram.memory\[138\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[0\]_D io_in[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08535__A1 _03547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07338__A2 _03255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10983_ _10983_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__10048__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05879__I u_cpu.cpu.bufreg.lsb\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10198__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09263__A2 _04506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05824__A2 u_cpu.cpu.bufreg.i_sh_signed vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09015__A2 _04369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05380__S0 _01546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10417_ _00850_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07577__A2 _03392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[19\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10348_ _00781_ io_in[4] u_cpu.rf_ram.memory\[121\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05588__A1 _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10279_ _00712_ io_in[4] u_cpu.rf_ram.memory\[91\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08526__A1 _02612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05119__I _01548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07329__A2 _03255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05563__B _01565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04840_ _01367_ _01368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_94_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05760__A1 _01609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06510_ u_cpu.rf_ram.memory\[16\]\[5\] _02791_ _02797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07490_ _03347_ _03345_ _03348_ _00624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07888__I0 _02587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05199__S0 _01687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07501__A2 _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06441_ _02748_ _02740_ _02749_ _00174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09160_ _04284_ _04449_ _04451_ _01192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06372_ u_cpu.rf_ram.memory\[43\]\[0\] _02708_ _02709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09833__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09254__A2 _04506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08111_ u_arbiter.i_wb_cpu_dbus_dat\[29\] _03723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06068__A2 _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05323_ u_cpu.rf_ram.memory\[36\]\[2\] u_cpu.rf_ram.memory\[37\]\[2\] u_cpu.rf_ram.memory\[38\]\[2\]
+ u_cpu.rf_ram.memory\[39\]\[2\] _01619_ _01620_ _01813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09091_ u_cpu.rf_ram.memory\[105\]\[3\] _04409_ _04413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08042_ _03654_ _03678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10810__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05254_ _01645_ _01744_ _01648_ _01745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_31_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09006__A2 _04359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05371__S0 _01680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07017__A1 _02957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09983__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05185_ _01670_ _01672_ _01674_ _01676_ _01568_ _01677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_89_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07568__A2 _03392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08765__A1 _02469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05579__A1 _01636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09993_ _00000_ io_in[4] u_cpu.rf_ram.rdata\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06240__A2 _02628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08944_ _04332_ _01095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08517__A1 _04016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08875_ u_cpu.rf_ram.memory\[94\]\[5\] _04282_ _04293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09190__A1 _04296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07826_ _03543_ _03541_ _03544_ _00765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07757_ u_cpu.rf_ram.memory\[92\]\[4\] _03500_ _03505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04969_ u_cpu.cpu.ctrl.o_ibus_adr\[12\] _01476_ u_cpu.cpu.ctrl.o_ibus_adr\[13\] _01480_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_25_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05751__A1 _01589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06708_ _02746_ _02904_ _02908_ _00282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07688_ _03462_ _00708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09493__A2 _04644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10340__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09427_ u_cpu.rf_ram.memory\[26\]\[4\] _04605_ _04610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06639_ u_cpu.rf_ram.memory\[74\]\[5\] _02864_ _02870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09358_ u_cpu.rf_ram.memory\[88\]\[7\] _04556_ _04564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_u_scanchain_local.scan_flop\[42\]_D u_scanchain_local.module_data_in\[41\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04857__A3 u_cpu.cpu.decode.op21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08309_ u_arbiter.i_wb_cpu_rdt\[5\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[5\]
+ _01436_ _03890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09289_ _04525_ _04526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10490__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05362__S0 _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07559__A2 _03382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10202_ _00648_ io_in[4] u_cpu.rf_ram.memory\[126\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10133_ _00579_ io_in[4] u_cpu.rf_ram.memory\[134\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08359__I1 u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10064_ _00510_ io_in[4] u_cpu.rf_ram.memory\[70\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05990__A1 _01387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[6\] u_arbiter.i_wb_cpu_rdt\[3\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[0\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__09706__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05383__B _01417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07731__A2 _03458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05742__A1 _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10966_ _10966_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__09856__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06298__A2 _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08692__B1 _04175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10897_ _01326_ io_in[4] u_cpu.rf_ram.memory\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10833__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[33\]_D u_arbiter.i_wb_cpu_rdt\[30\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07798__A2 _03520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05353__S0 _01590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06470__A2 u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08747__A1 _03555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06222__A2 _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10213__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06990_ u_cpu.rf_ram.memory\[55\]\[6\] _03061_ _03068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05941_ _02321_ u_cpu.rf_ram.rdata\[4\] _02418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09172__A1 _04296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08660_ u_arbiter.i_wb_cpu_ibus_adr\[1\] _04155_ _04157_ u_cpu.cpu.ctrl.o_ibus_adr\[2\]
+ _04159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05872_ _01370_ _02351_ _02353_ _02354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_54_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07722__A2 _03475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09480__S _04634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07611_ u_cpu.rf_ram.memory\[123\]\[5\] _03412_ _03418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10363__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08591_ u_arbiter.i_wb_cpu_dbus_adr\[16\] u_arbiter.i_wb_cpu_dbus_adr\[15\] _04115_
+ _04118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__05733__A1 _01542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07542_ _03357_ _03372_ _03379_ _00645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06289__A2 _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07473_ _02587_ u_cpu.rf_ram.memory\[12\]\[3\] _03334_ _03338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_35_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07486__A1 u_cpu.rf_ram.memory\[22\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05740__C _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09212_ u_cpu.rf_ram.memory\[84\]\[6\] _04470_ _04483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06424_ _02517_ _02729_ _02737_ _00169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[24\]_D u_arbiter.i_wb_cpu_rdt\[21\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09227__A2 _04487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07238__A1 _03161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06355_ u_cpu.rf_ram.memory\[41\]\[1\] _02697_ _02699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09143_ u_cpu.rf_ram.memory\[83\]\[2\] _04439_ _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07789__A2 _03520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08986__A1 _04290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05306_ _01570_ _01795_ _01796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09074_ _04288_ _04399_ _04403_ _01154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06286_ _02507_ _02651_ _02657_ _00111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05237_ u_cpu.rf_ram.memory\[32\]\[1\] u_cpu.rf_ram.memory\[33\]\[1\] u_cpu.rf_ram.memory\[34\]\[1\]
+ u_cpu.rf_ram.memory\[35\]\[1\] _01623_ _01624_ _01728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_107_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08025_ u_arbiter.i_wb_cpu_dbus_dat\[0\] u_arbiter.i_wb_cpu_dbus_dat\[1\] u_arbiter.i_wb_cpu_dbus_dat\[2\]
+ _02774_ _03663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_104_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05168_ u_cpu.rf_ram.memory\[88\]\[0\] u_cpu.rf_ram.memory\[89\]\[0\] u_cpu.rf_ram.memory\[90\]\[0\]
+ u_cpu.rf_ram.memory\[91\]\[0\] _01646_ _01624_ _01660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_104_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09729__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09976_ _00430_ io_in[4] u_cpu.rf_ram.memory\[52\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05099_ _01548_ _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07961__A2 _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08927_ _04280_ _04322_ _04323_ _01087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10706__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05972__A1 _01374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08858_ _02475_ _02625_ _04281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09879__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07713__A2 _03475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08910__A1 _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07903__S _03586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07809_ u_cpu.rf_ram.memory\[117\]\[3\] _03530_ _03534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05724__A1 _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08789_ _03545_ _04227_ _04230_ _01042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10820_ _01249_ io_in[4] u_cpu.rf_ram.memory\[86\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10856__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09466__A2 _04625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10751_ _01180_ io_in[4] u_cpu.rf_ram.memory\[107\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08674__B1 _04157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[15\]_D u_arbiter.i_wb_cpu_rdt\[12\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10682_ _01111_ io_in[4] u_cpu.rf_ram.memory\[101\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05583__S0 _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08277__I0 u_arbiter.i_wb_cpu_rdt\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10236__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08729__A1 u_cpu.cpu.immdec.imm11_7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07401__A1 _03163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10116_ _00562_ io_in[4] u_cpu.rf_ram.memory\[136\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10386__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11096_ _11096_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_95_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05963__A1 _01403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09154__A1 _04296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10047_ _00493_ io_in[4] u_cpu.rf_ram.memory\[73\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07704__A2 _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08901__A1 _02612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05715__A1 _01667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05191__A2 _01682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09457__A2 _04625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10949_ u_cpu.rf_ram_if.wdata1_r\[3\] io_in[4] u_cpu.rf_ram_if.wdata1_r\[2\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09209__A2 _04470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06140__A1 _02482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05132__I _01547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05574__S0 _01590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06140_ _02482_ _02563_ _02564_ _00058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06164__S _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08432__A3 _03770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07640__A1 _03347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06071_ _01547_ _02519_ _02520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__05288__B _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06443__A2 _02740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05022_ u_cpu.cpu.ctrl.o_ibus_adr\[25\] u_cpu.cpu.ctrl.o_ibus_adr\[24\] _01513_ _01520_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_113_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10729__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08196__A2 u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09830_ _00284_ io_in[4] u_cpu.rf_ram.memory\[68\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07943__A2 _03606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09761_ _00215_ io_in[4] u_cpu.rf_ram.memory\[119\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06973_ _02967_ _03051_ _03058_ _00397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08712_ u_cpu.cpu.ctrl.o_ibus_adr\[26\] _04173_ _04175_ u_cpu.cpu.ctrl.o_ibus_adr\[27\]
+ _04186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_132_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05924_ _02403_ _02398_ _02399_ _02405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_09692_ _00146_ io_in[4] u_cpu.rf_ram.memory\[43\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10879__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08643_ _03545_ _04145_ _04148_ _00978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05706__A1 _01609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05855_ u_cpu.cpu.mem_bytecnt\[1\] u_cpu.cpu.state.o_cnt\[2\] u_cpu.cpu.mem_bytecnt\[0\]
+ _02338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_82_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08574_ u_arbiter.i_wb_cpu_dbus_adr\[8\] u_arbiter.i_wb_cpu_dbus_adr\[7\] _02445_
+ _04109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05786_ _01614_ _02270_ _01626_ _02271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09448__A2 _04615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05182__A2 _01673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10109__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07459__A1 _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07525_ u_cpu.rf_ram.memory\[128\]\[7\] _03362_ _03370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08120__A2 _02781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07456_ u_cpu.rf_ram.memory\[130\]\[3\] _03325_ _03329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05565__S0 _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06407_ _02639_ _02727_ _02728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06682__A2 _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10259__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07387_ _03167_ _03285_ _03290_ _00579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09126_ _04286_ _04429_ _04432_ _01177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06338_ u_cpu.rf_ram.memory\[51\]\[2\] _02686_ _02689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09057_ u_cpu.rf_ram.memory\[99\]\[4\] _04389_ _04394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06269_ u_cpu.rf_ram.memory\[42\]\[6\] _02641_ _02648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06434__A2 _02740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08008_ _02772_ _03647_ _03648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08187__A2 _03778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09959_ _00413_ io_in[4] u_cpu.rf_ram.memory\[54\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05945__A1 _02320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09136__A1 _04296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06370__A1 _02639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05173__A2 _01664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09439__A2 _04615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10803_ _01232_ io_in[4] u_cpu.rf_ram.memory\[85\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08498__I0 u_arbiter.i_wb_cpu_rdt\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10734_ _01163_ io_in[4] u_cpu.rf_ram.memory\[105\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06122__A1 _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05556__S0 _01546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07870__A1 _03545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06673__A2 _02884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10665_ _01094_ io_in[4] u_cpu.rf_ram.memory\[28\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10596_ _01025_ io_in[4] u_cpu.rf_ram.memory\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07622__A1 _03347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[43\] u_scanchain_local.module_data_in\[42\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[5\] u_scanchain_local.clk u_scanchain_local.module_data_in\[43\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04987__A2 _01457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08178__A2 u_arbiter.i_wb_cpu_rdt\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09375__A1 _04568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07925__A2 _03596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05936__A1 _02320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11079_ _11079_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_110_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05127__I _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07689__A1 _01428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08350__A2 _03768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05640_ _01684_ _02126_ _01418_ _02127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_91_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05795__S0 _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05571_ u_cpu.rf_ram.memory\[24\]\[5\] u_cpu.rf_ram.memory\[25\]\[5\] u_cpu.rf_ram.memory\[26\]\[5\]
+ u_cpu.rf_ram.memory\[27\]\[5\] _01578_ _01580_ _02058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_16_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07310_ u_cpu.rf_ram.memory\[137\]\[2\] _03245_ _03248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10401__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08290_ _03878_ _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05547__S0 _01680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09574__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07241_ u_cpu.rf_ram.memory\[143\]\[3\] _03206_ _03210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07172_ _03169_ _03159_ _03170_ _00484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06123_ u_cpu.rf_ram.memory\[18\]\[2\] _02551_ _02554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10551__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06416__A2 _02729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06054_ _02505_ _02506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04978__A2 u_cpu.cpu.ctrl.o_ibus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08169__A2 _03768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05005_ u_cpu.cpu.ctrl.o_ibus_adr\[21\] u_cpu.cpu.ctrl.o_ibus_adr\[20\] u_cpu.cpu.ctrl.o_ibus_adr\[19\]
+ _01495_ _01507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_99_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09813_ _00267_ io_in[4] u_cpu.rf_ram.memory\[75\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05465__C _01404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09118__A1 _04296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09744_ _00198_ io_in[4] u_cpu.rf_ram.memory\[16\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_101_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06956_ u_cpu.rf_ram.memory\[57\]\[7\] _03041_ _03049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05907_ _01369_ _02387_ _02388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09675_ _00129_ io_in[4] u_cpu.rf_ram.memory\[44\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06887_ _02528_ _02682_ _03011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08341__A2 _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08626_ _02444_ _02773_ _04136_ _04137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_43_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05838_ u_cpu.rf_ram.rdata\[0\] _02321_ _02322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08557_ _03551_ _04094_ _04100_ _00940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09917__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05769_ _01539_ _02225_ _02234_ _02253_ _02254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_70_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10081__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07508_ _03359_ _03345_ _03360_ _00630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06104__A1 _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05538__S0 _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08488_ u_arbiter.i_wb_cpu_rdt\[17\] u_arbiter.i_wb_cpu_rdt\[1\] _01436_ _04050_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_74_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07852__A1 _03545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06655__A2 _02874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07439_ _03165_ _03315_ _03319_ _00602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10450_ _00883_ io_in[4] u_cpu.rf_ram.memory\[113\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09109_ u_cpu.rf_ram.memory\[106\]\[3\] _04419_ _04423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07604__A1 _03347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06407__A2 _02727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10381_ _00814_ io_in[4] u_cpu.rf_ram.memory\[122\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05710__S0 _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05091__A1 _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09357__A1 _04482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05656__B _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11002_ _11002_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_105_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[52\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05918__A1 _02361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06591__A1 _02706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[12\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10424__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06343__A1 _02502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09597__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06894__A2 _03012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[27\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08096__A1 u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05529__S0 _01590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07143__I0 _02587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10574__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10717_ _01146_ io_in[4] u_cpu.rf_ram.memory\[99\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10648_ _01077_ io_in[4] u_cpu.rf_ram.memory\[96\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10579_ _01009_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05701__S0 _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08020__A1 u_arbiter.i_wb_cpu_dbus_dat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05909__A1 _02381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06810_ u_cpu.rf_ram.memory\[29\]\[6\] _02955_ _02968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07790_ _03349_ _03520_ _03523_ _00750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05385__A2 _01873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06582__A1 _02746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06741_ u_cpu.rf_ram.memory\[66\]\[2\] _02924_ _02927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09460_ _04474_ _04625_ _04628_ _01315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05137__A2 _01618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06672_ _02746_ _02884_ _02888_ _00266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08411_ _03897_ _03981_ _03906_ _03982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_24_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05623_ _01667_ _02109_ _02110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10917__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09391_ u_cpu.cpu.genblk3.csr.mstatus_mpie _01377_ _01393_ _04589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06885__A2 _03002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08342_ _03866_ _03920_ _00905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05554_ _02032_ _02041_ _02042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06637__A2 _02864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08273_ _03800_ _03859_ _03863_ _03761_ _03864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05485_ _01966_ _01968_ _01970_ _01972_ _01426_ _01973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_07224_ _03165_ _03196_ _03200_ _00506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07155_ _03158_ _03159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06106_ _02492_ _02541_ _02544_ _00044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07086_ u_cpu.rf_ram.memory\[142\]\[1\] _03119_ _03121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09339__A1 _04482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06037_ _02491_ _02492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05612__A3 _02098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08011__A1 u_arbiter.i_wb_cpu_dbus_dat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08562__A2 _02433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10447__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07988_ _03635_ _03636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05376__A2 _01865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06573__A1 _02539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09727_ _00181_ io_in[4] u_cpu.rf_ram.memory\[4\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06939_ _02969_ _03031_ _03039_ _00382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09511__A1 _04472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09658_ _00112_ io_in[4] u_cpu.rf_ram.memory\[46\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05759__S0 _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07911__S _03586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10597__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08609_ u_arbiter.i_wb_cpu_dbus_adr\[25\] u_arbiter.i_wb_cpu_dbus_adr\[24\] _04115_
+ _04127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_76_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06876__A2 _03002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09589_ _00043_ io_in[4] u_cpu.rf_ram.memory\[81\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__04887__A1 _01411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08078__A1 u_arbiter.i_wb_cpu_rdt\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08078__B2 u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10502_ _00935_ io_in[4] u_cpu.rf_ram.memory\[31\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10433_ _00866_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08250__A1 _03762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10364_ _00797_ io_in[4] u_cpu.rf_ram.memory\[11\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10295_ _00728_ io_in[4] u_cpu.cpu.mem_if.signbit vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08002__A1 _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06061__I _02511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08553__A2 _04094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05367__A2 _01847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08305__A2 _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06316__A1 _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06867__A2 _02992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__04878__A1 _01377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08069__A1 u_arbiter.i_wb_cpu_dbus_dat\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07816__A1 _03357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06619__A2 _02854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05270_ u_cpu.rf_ram.memory\[64\]\[1\] u_cpu.rf_ram.memory\[65\]\[1\] u_cpu.rf_ram.memory\[66\]\[1\]
+ u_cpu.rf_ram.memory\[67\]\[1\] _01571_ _01668_ _01761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07292__A2 _03235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09612__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08241__A1 _03751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06172__S _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07044__A2 _03091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08792__A2 _04227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08960_ _04340_ _01103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07911_ _02596_ u_cpu.rf_ram.memory\[11\]\[6\] _03586_ _03593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_111_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08891_ u_cpu.rf_ram.memory\[95\]\[3\] _04299_ _04303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09762__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08544__A2 _02727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07842_ _02516_ _03555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07773_ u_cpu.rf_ram.memory\[35\]\[3\] _03510_ _03514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04985_ _01443_ _01490_ _01491_ _01492_ u_arbiter.o_wb_cpu_adr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_09512_ u_cpu.rf_ram.memory\[100\]\[2\] _04654_ _04657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06724_ _02744_ _02914_ _02917_ _00289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06307__A1 _02512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09443_ u_cpu.rf_ram.memory\[25\]\[3\] _04615_ _04619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06655_ u_cpu.rf_ram.memory\[76\]\[4\] _02874_ _02879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06858__A2 _02992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__04869__A1 _01393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05606_ _01601_ _02092_ _01648_ _02093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_12_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09374_ u_cpu.cpu.genblk3.csr.mcause3_0\[2\] _04568_ _04577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06586_ _02750_ _02834_ _02840_ _00228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08325_ _03831_ _03897_ _03791_ _03906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05537_ _01553_ _02024_ _01565_ _02025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_138_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08256_ _03763_ _03785_ _03809_ _03848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07283__A2 _03225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05468_ u_cpu.rf_ram.memory\[8\]\[4\] u_cpu.rf_ram.memory\[9\]\[4\] u_cpu.rf_ram.memory\[10\]\[4\]
+ u_cpu.rf_ram.memory\[11\]\[4\] _01546_ _01550_ _01956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__05050__I _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07207_ u_cpu.rf_ram.memory\[71\]\[4\] _03186_ _03191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08187_ _03776_ _03778_ _03787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05833__A3 _01374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05399_ _01589_ _01887_ _01888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08232__A1 _03757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07138_ _03149_ _00471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07035__A2 _03091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07069_ _03111_ _00440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_79_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05597__A2 _02083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10080_ _00526_ io_in[4] u_cpu.rf_ram.memory\[14\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08535__A2 _04084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06546__A1 _02748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10982_ _10982_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_74_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06849__A2 _02982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09635__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08471__A1 _03768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07274__A2 _03225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05904__S0 u_cpu.cpu.bufreg.lsb\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05675__I3 u_cpu.rf_ram.memory\[39\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05380__S1 _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10612__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10416_ _00849_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08223__A1 _03818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07026__A2 _03081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05037__A1 _01443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09785__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10347_ _00780_ io_in[4] u_cpu.rf_ram.memory\[121\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10278_ _00711_ io_in[4] u_cpu.rf_ram.memory\[91\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10762__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08526__A2 _02639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[5\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05760__A2 _02244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05199__S1 _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06440_ u_cpu.rf_ram.memory\[50\]\[4\] _02740_ _02749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10142__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06371_ _02707_ _02708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09478__S _04634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08110_ _03721_ _03722_ _00871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05322_ _01614_ _01811_ _01605_ _01812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09090_ _04286_ _04409_ _04412_ _01161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08462__A1 _03751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08041_ u_arbiter.i_wb_cpu_dbus_dat\[5\] _02774_ _03674_ _03676_ _03677_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05253_ u_cpu.rf_ram.memory\[120\]\[1\] u_cpu.rf_ram.memory\[121\]\[1\] u_cpu.rf_ram.memory\[122\]\[1\]
+ u_cpu.rf_ram.memory\[123\]\[1\] _01646_ _01603_ _01744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10292__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05371__S1 _01681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08214__A1 _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07017__A2 _03081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05184_ _01636_ _01675_ _01417_ _01676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08765__A2 _02577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09992_ _00446_ io_in[4] u_cpu.rf_ram.memory\[15\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05579__A2 _02065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06776__A1 _02742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08943_ u_arbiter.i_wb_cpu_rdt\[16\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[0\]
+ _04331_ _04332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08874_ _02506_ _04292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07825_ u_cpu.rf_ram.memory\[120\]\[1\] _03541_ _03544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09190__A2 _04459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05200__A1 _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07756_ _03351_ _03500_ _03504_ _00735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04968_ _01445_ _01478_ _01479_ u_arbiter.o_wb_cpu_adr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06707_ u_cpu.rf_ram.memory\[68\]\[3\] _02904_ _02908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07687_ _01429_ u_cpu.cpu.state.o_cnt_r\[0\] _03462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_04899_ _01423_ _01424_ _01425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09426_ _04476_ _04605_ _04609_ _01300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09658__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06638_ _02748_ _02864_ _02869_ _00251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_125_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09357_ _04482_ _04556_ _04563_ _01277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06569_ _02752_ _02823_ _02830_ _00221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__04857__A4 u_cpu.cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10635__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08308_ _03816_ _03888_ _03889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09288_ _02475_ _02893_ _04525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08453__B2 _03834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08239_ _03740_ _03833_ _03834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05362__S1 _01668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08205__A1 _03801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07008__A2 _03071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10785__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10201_ _00647_ io_in[4] u_cpu.rf_ram.memory\[126\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10132_ _00578_ io_in[4] u_cpu.rf_ram.memory\[134\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10015__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10063_ _00509_ io_in[4] u_cpu.rf_ram.memory\[70\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06519__A1 _02738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05990__A2 _02433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09181__A2 _04459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07192__A1 _03169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10165__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10965_ _10965_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_62_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07495__A2 _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10896_ _01325_ io_in[4] u_cpu.rf_ram.memory\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07170__I _02506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08444__A1 _04010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07247__A2 _03206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08444__B2 _03798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05258__A1 _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08995__A2 _04359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05353__S1 _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08215__B _03812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09244__I0 _02590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08747__A2 _04199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06758__A1 _02742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05430__A1 _01645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05940_ _02320_ _02416_ _02417_ _00017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_65_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09172__A2 _04449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05871_ u_cpu.cpu.bne_or_bge _02351_ _02352_ _02353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10508__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07610_ _03353_ _03412_ _03417_ _00675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08590_ _04117_ _00956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09800__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05733__A2 _02217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07541_ u_cpu.rf_ram.memory\[127\]\[6\] _03372_ _03379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10658__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07472_ _03337_ _00617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07486__A2 _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09211_ _02511_ _04482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06423_ u_cpu.rf_ram.memory\[47\]\[7\] _02729_ _02737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09950__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09142_ _04284_ _04439_ _04441_ _01184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06354_ _02482_ _02697_ _02698_ _00138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08435__A1 _03999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07238__A2 _03206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05249__A1 _01601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05305_ u_cpu.rf_ram.memory\[28\]\[2\] u_cpu.rf_ram.memory\[29\]\[2\] u_cpu.rf_ram.memory\[30\]\[2\]
+ u_cpu.rf_ram.memory\[31\]\[2\] _01572_ _01574_ _01795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08986__A2 _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09073_ u_cpu.rf_ram.memory\[79\]\[3\] _04399_ _04403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06285_ u_cpu.rf_ram.memory\[46\]\[5\] _02651_ _02657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06997__A1 _02953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08024_ u_arbiter.i_wb_cpu_dbus_dat\[3\] _02774_ _03662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05236_ _01589_ _01726_ _01727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08738__A2 _04199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10038__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05167_ _01398_ _01658_ _01659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05098_ _01544_ _01590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09975_ _00429_ io_in[4] u_cpu.rf_ram.memory\[52\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07410__A2 _03295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05421__A1 _01594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08926_ u_cpu.rf_ram.memory\[28\]\[0\] _04322_ _04323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05484__B _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05972__A2 u_cpu.cpu.decode.opcode\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09163__A2 _04449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10188__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08857_ _02481_ _04280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08910__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07808_ _03349_ _03530_ _03533_ _00758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08788_ u_cpu.rf_ram.memory\[93\]\[2\] _04227_ _04230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05724__A2 _02209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[3\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07739_ _03491_ _03492_ _03493_ _02359_ _03494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_77_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10750_ _01179_ io_in[4] u_cpu.rf_ram.memory\[107\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09409_ u_cpu.rf_ram.memory\[27\]\[4\] _04595_ _04600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10681_ _01110_ io_in[4] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05583__S1 _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07229__A2 _03196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08277__I1 u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09474__I0 _02581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08977__A2 _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08035__B _03653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05660__A1 _01542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07401__A2 _03295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05412__A1 _01589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06460__I0 _02590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10115_ _00561_ io_in[4] u_cpu.rf_ram.memory\[136\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11095_ _11095_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_1_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09823__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09154__A2 _04439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10046_ _00492_ io_in[4] u_cpu.rf_ram.memory\[73\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08901__A2 _04197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05715__A2 _02200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10800__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09973__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10948_ u_cpu.rf_ram_if.wdata1_r\[2\] io_in[4] u_cpu.rf_ram_if.wdata1_r\[1\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10879_ _01308_ io_in[4] u_cpu.rf_ram.memory\[25\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10950__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06140__A2 _02563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05574__S1 _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08417__A1 _03741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09090__A1 _04286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06979__A1 _02953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06070_ u_cpu.rf_ram_if.rcnt\[1\] u_cpu.rf_ram_if.rcnt\[0\] _01543_ u_cpu.rf_ram_if.rcnt\[2\]
+ _02519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__07640__A2 _03432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05651__A1 _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05021_ _01445_ _01518_ _01519_ u_arbiter.o_wb_cpu_adr\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06180__S _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10330__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05403__A1 _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09760_ _00214_ io_in[4] u_cpu.rf_ram.memory\[40\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06972_ u_cpu.rf_ram.memory\[56\]\[6\] _03051_ _03058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05954__A2 _01403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08711_ _04185_ _01009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__09145__A2 _04439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05923_ _02398_ _02399_ _02403_ _02404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09691_ _00145_ io_in[4] u_cpu.rf_ram.memory\[41\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06203__I0 _02590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08642_ u_cpu.rf_ram.memory\[30\]\[2\] _04145_ _04148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10480__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05854_ u_cpu.cpu.decode.op22 _02337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_39_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05706__A2 _02191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08573_ _04108_ _00948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05785_ u_cpu.rf_ram.memory\[116\]\[7\] u_cpu.rf_ram.memory\[117\]\[7\] u_cpu.rf_ram.memory\[118\]\[7\]
+ u_cpu.rf_ram.memory\[119\]\[7\] _01623_ _01624_ _02270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_42_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07524_ _03357_ _03362_ _03369_ _00637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08656__A1 _01428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07459__A2 _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07455_ _03163_ _03325_ _03328_ _00609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06131__A2 _02551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05565__S1 _01574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06406_ _02601_ _02624_ _02727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_10_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08408__A1 _02765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07386_ u_cpu.rf_ram.memory\[134\]\[4\] _03285_ _03290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09125_ u_cpu.rf_ram.memory\[107\]\[2\] _04429_ _04432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06337_ _02487_ _02686_ _02688_ _00131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09056_ _04288_ _04389_ _04393_ _01146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07631__A2 _03422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06268_ _02507_ _02641_ _02647_ _00103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08570__S _02445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08007_ _02305_ _03645_ _03646_ _03647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__05642__A1 _02119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05219_ u_cpu.rf_ram.memory\[24\]\[1\] u_cpu.rf_ram.memory\[25\]\[1\] u_cpu.rf_ram.memory\[26\]\[1\]
+ u_cpu.rf_ram.memory\[27\]\[1\] _01578_ _01580_ _01710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_144_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06199_ _02584_ u_cpu.rf_ram.memory\[7\]\[2\] _02603_ _02606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09846__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09958_ _00412_ io_in[4] u_cpu.rf_ram.memory\[54\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10823__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09136__A2 _04429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08909_ u_cpu.rf_ram.memory\[96\]\[3\] _04309_ _04313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09889_ _00343_ io_in[4] u_cpu.rf_ram.memory\[61\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09996__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07698__A2 _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05253__S0 _01646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05661__C _01426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06370__A2 _02706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10802_ _01231_ io_in[4] u_cpu.rf_ram.memory\[85\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08647__A1 _03549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08498__I1 u_arbiter.i_wb_cpu_rdt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10733_ _01162_ io_in[4] u_cpu.rf_ram.memory\[105\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06122__A2 _02551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05556__S1 _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10203__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10664_ _01093_ io_in[4] u_cpu.rf_ram.memory\[28\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07870__A2 _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09072__A1 _04286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10595_ _01024_ io_in[4] u_cpu.rf_ram.memory\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07622__A2 _03422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10353__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_scanchain_local.scan_flop\[36\] u_scanchain_local.module_data_in\[35\] io_in[3]
+ u_arbiter.i_wb_cpu_dbus_dat\[30\] u_scanchain_local.clk u_scanchain_local.module_data_in\[36\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_135_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09127__A2 _04429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05492__S0 _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11078_ _11078_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_62_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05852__B _02333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10029_ _00475_ io_in[4] u_cpu.rf_ram.memory\[13\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05149__B1 _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08886__A1 _04280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05244__S0 _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06361__A2 _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05795__S1 _01652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05570_ _01570_ _02056_ _02057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09719__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06113__A2 _02541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05547__S1 _01681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07240_ _03163_ _03206_ _03209_ _00513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07861__A2 _03558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05872__A1 _01370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07171_ u_cpu.rf_ram.memory\[72\]\[5\] _03159_ _03170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05299__B _01565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09486__S _04634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09869__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06122_ _02487_ _02551_ _02553_ _00051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08390__S _01437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07613__A2 _03412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08810__A1 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06053_ _02460_ u_cpu.rf_ram_if.wdata0_r\[5\] _02504_ _02505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10846__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05004_ u_cpu.cpu.ctrl.o_ibus_adr\[22\] _01506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_28_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09812_ _00266_ io_in[4] u_cpu.rf_ram.memory\[75\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09118__A2 _04419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05483__S0 _01578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06955_ _02967_ _03041_ _03048_ _00389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09743_ _00197_ io_in[4] u_cpu.rf_ram.memory\[16\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07129__A1 _02963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05762__B _01416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05906_ _02384_ _02385_ _02387_ _00728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09674_ _00128_ io_in[4] u_cpu.rf_ram.memory\[44\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06886_ _02969_ _03002_ _03010_ _00358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05235__S0 _01619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08625_ _01372_ _02394_ _02441_ _02443_ _04136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_43_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05837_ u_cpu.rf_ram.regzero _02321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_82_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10226__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08629__A1 _02372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08556_ u_cpu.rf_ram.memory\[31\]\[5\] _04094_ _04100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05768_ _01421_ _02243_ _02252_ _02253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__05053__I _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07507_ u_cpu.rf_ram.memory\[22\]\[7\] _03345_ _03360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08487_ _04016_ _04047_ _04048_ _04049_ _00921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_126_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05699_ _02178_ _02180_ _02182_ _02184_ _01607_ _02185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__06104__A2 _02541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07301__A1 _03171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05538__S1 _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04892__I _01417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07438_ u_cpu.rf_ram.memory\[131\]\[3\] _03315_ _03319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07852__A2 _03558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10376__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05863__A1 _02341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09054__A1 _04286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07369_ _03167_ _03275_ _03280_ _00571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09108_ _04286_ _04419_ _04422_ _01169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07909__S _03586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07604__A2 _03412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10380_ _00813_ io_in[4] u_cpu.rf_ram.memory\[122\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08801__A1 _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09039_ u_cpu.rf_ram.memory\[104\]\[4\] _04379_ _04384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05710__S1 _01668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09357__A2 _04556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05091__A2 _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11001_ _11001_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_104_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06040__A1 _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09109__A2 _04419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05474__S0 _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08168__I0 u_arbiter.i_wb_cpu_rdt\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06591__A2 _02832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05226__S0 _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07540__A1 _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06343__A2 _02686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10719__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09293__A1 _04472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08096__A2 _03683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05529__S1 _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10716_ _01145_ io_in[4] u_cpu.rf_ram.memory\[99\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07843__A2 _03541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10647_ _01076_ io_in[4] u_cpu.rf_ram.memory\[95\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10869__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10578_ _01008_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05606__A1 _01601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05701__S1 _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08223__B _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09348__A2 _04556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06582__A2 _02834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10249__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06740_ _02742_ _02924_ _02926_ _00296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05217__S0 _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09520__A2 _04654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06671_ u_cpu.rf_ram.memory\[75\]\[3\] _02884_ _02888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06334__A2 _02686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08410_ _03742_ _03786_ _03902_ _03899_ _03981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_52_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05622_ u_cpu.rf_ram.memory\[64\]\[5\] u_cpu.rf_ram.memory\[65\]\[5\] u_cpu.rf_ram.memory\[66\]\[5\]
+ u_cpu.rf_ram.memory\[67\]\[5\] _01571_ _01668_ _02109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09390_ _04191_ _02348_ _04588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10399__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08341_ u_cpu.cpu.immdec.imm24_20\[1\] _03916_ _03919_ u_cpu.cpu.immdec.imm24_20\[2\]
+ _03920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05553_ _02034_ _02036_ _02038_ _02040_ _01404_ _02041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_71_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09691__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08272_ _03773_ _03860_ _03862_ _03755_ _03863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__07834__A2 _03541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05484_ _01542_ _01971_ _01418_ _01972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07223_ u_cpu.rf_ram.memory\[70\]\[3\] _03196_ _03200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05845__A1 _02305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09036__A1 _04286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07154_ _02626_ _02810_ _03158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07598__A1 _03359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06105_ u_cpu.rf_ram.memory\[81\]\[2\] _02541_ _02544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05757__B _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07085_ _02953_ _03119_ _03120_ _00447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06270__A1 _02512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09339__A2 _04546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06036_ _02490_ _02491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05476__C _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08011__A2 _02774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07070__I0 _02584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07987_ _02539_ _02639_ _03635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07770__A1 _03347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06573__A2 _02832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09726_ _00180_ io_in[4] u_cpu.rf_ram.memory\[4\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06938_ u_cpu.rf_ram.memory\[58\]\[7\] _03031_ _03039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05208__S0 _01546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09511__A2 _04654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09657_ _00111_ io_in[4] u_cpu.rf_ram.memory\[46\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06869_ _02671_ _02684_ _03001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06325__A2 _02673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07522__A1 _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05759__S1 _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08608_ _04126_ _00965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_70_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09588_ _00042_ io_in[4] u_cpu.rf_ram.memory\[81\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08539_ _03551_ _04084_ _04090_ _00932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04887__A2 _01412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09275__A1 _04472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08078__A2 _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06089__A1 _02497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07825__A2 _03541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10501_ _00934_ io_in[4] u_cpu.rf_ram.memory\[32\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10432_ _00865_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10363_ _00796_ io_in[4] u_cpu.rf_ram.memory\[11\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08250__A2 _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05695__S0 _01619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10294_ _00727_ io_in[4] u_cpu.cpu.state.genblk1.misalign_trap_sync_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08002__A2 _03636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06013__A1 u_cpu.cpu.immdec.imm11_7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07061__I0 _02596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06564__A2 _02823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05367__A3 _01856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07173__I _02511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09502__A2 _04644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10541__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06316__A2 _02673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08710__B1 _04175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__04878__A2 _01387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08069__A2 _03683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10691__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07816__A2 _03530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09018__A1 _04286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05577__B _01564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05686__S0 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07910_ _03592_ _00801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09907__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08890_ _04286_ _04299_ _04302_ _01071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10071__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07841_ _03553_ _03541_ _03554_ _00770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07752__A1 _03347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07772_ _03349_ _03510_ _03513_ _00742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_04984_ u_arbiter.i_wb_cpu_dbus_adr\[16\] _01442_ _01492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09511_ _04472_ _04654_ _04656_ _01338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06723_ u_cpu.rf_ram.memory\[67\]\[2\] _02914_ _02917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06307__A2 _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07504__A1 u_cpu.rf_ram.memory\[22\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09442_ _04474_ _04615_ _04618_ _01307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06654_ _02746_ _02874_ _02878_ _00258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05605_ u_cpu.rf_ram.memory\[120\]\[5\] u_cpu.rf_ram.memory\[121\]\[5\] u_cpu.rf_ram.memory\[122\]\[5\]
+ u_cpu.rf_ram.memory\[123\]\[5\] _01646_ _01603_ _02092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04869__A2 _01394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09373_ u_cpu.cpu.genblk3.csr.mcause3_0\[3\] _01393_ u_cpu.cpu.genblk3.csr.o_new_irq
+ _01375_ _04576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__09257__A1 _04472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06585_ u_cpu.rf_ram.memory\[129\]\[5\] _02834_ _02840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08324_ _03744_ _03786_ _03828_ _03890_ _03904_ _03905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_05536_ u_cpu.rf_ram.memory\[68\]\[4\] u_cpu.rf_ram.memory\[69\]\[4\] u_cpu.rf_ram.memory\[70\]\[4\]
+ u_cpu.rf_ram.memory\[71\]\[4\] _01555_ _01652_ _02024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07807__A2 _03530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[42\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05818__A1 _02293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08255_ _03752_ _03770_ _03787_ _03763_ _03800_ _03847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_05467_ _01406_ _01906_ _01955_ _00003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08480__A2 _04041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07206_ _03165_ _03186_ _03190_ _00498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08186_ _03776_ _03785_ _03786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08607__I1 u_arbiter.i_wb_cpu_dbus_adr\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05398_ u_cpu.rf_ram.memory\[52\]\[3\] u_cpu.rf_ram.memory\[53\]\[3\] u_cpu.rf_ram.memory\[54\]\[3\]
+ u_cpu.rf_ram.memory\[55\]\[3\] _01590_ _01591_ _01887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_4_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[11\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07137_ _02573_ u_cpu.rf_ram.memory\[13\]\[0\] _03148_ _03149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08232__A2 _03759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10414__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06243__A1 _02497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05677__S0 _01623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07068_ _02581_ u_cpu.rf_ram.memory\[15\]\[1\] _03109_ _03111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_134_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09587__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06019_ _02469_ _02475_ _02476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05841__I1 _02324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[26\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05429__S0 _01646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10564__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06546__A2 _02812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07743__A1 u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09709_ _00163_ io_in[4] u_cpu.rf_ram.memory\[47\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10981_ _10981_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__08299__A2 _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08753__S _04208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08471__A2 _03774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05904__S1 u_cpu.cpu.bufreg.lsb\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06482__A1 _02774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10415_ _00848_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09420__A1 _04468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10094__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06234__A1 _02625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10346_ _00779_ io_in[4] u_cpu.rf_ram.memory\[118\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05668__S0 _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07982__A1 _03551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06785__A2 _02944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10907__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10277_ _00710_ io_in[4] u_cpu.cpu.state.o_cnt_r\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06800__I _02496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06537__A2 _02812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07734__A1 _02325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[65\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06370_ _02639_ _02706_ _02707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05321_ u_cpu.rf_ram.memory\[44\]\[2\] u_cpu.rf_ram.memory\[45\]\[2\] u_cpu.rf_ram.memory\[46\]\[2\]
+ u_cpu.rf_ram.memory\[47\]\[2\] _01615_ _01616_ _01811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_30_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08462__A2 _03765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10437__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08040_ _03675_ _03676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06473__A1 _01428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05252_ _01398_ _01742_ _01743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05183_ u_cpu.rf_ram.memory\[76\]\[0\] u_cpu.rf_ram.memory\[77\]\[0\] u_cpu.rf_ram.memory\[78\]\[0\]
+ u_cpu.rf_ram.memory\[79\]\[0\] _01577_ _01549_ _01675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_31_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06225__A1 _02507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05028__A2 _01457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05659__S0 _01578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10587__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09991_ _00445_ io_in[4] u_cpu.rf_ram.memory\[15\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06776__A2 _02944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08942_ _02766_ _04331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08411__B _03906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08517__A3 _04075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08873_ _04290_ _04282_ _04291_ _01065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07725__A1 _03357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06528__A2 _02801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07824_ _02486_ _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05200__A2 _01691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07755_ u_cpu.rf_ram.memory\[92\]\[3\] _03500_ _03504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04967_ u_arbiter.i_wb_cpu_dbus_adr\[12\] _01457_ _01479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06706_ _02744_ _02904_ _02907_ _00281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07686_ _03459_ _03461_ _00707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04898_ u_cpu.cpu.immdec.imm24_20\[2\] _01388_ _01424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08150__A1 _01436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06637_ u_cpu.rf_ram.memory\[74\]\[4\] _02864_ _02869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09425_ u_cpu.rf_ram.memory\[26\]\[3\] _04605_ _04609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09356_ u_cpu.rf_ram.memory\[88\]\[6\] _04556_ _04563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06568_ u_cpu.rf_ram.memory\[119\]\[6\] _02823_ _02830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05061__I _01397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05519_ u_cpu.rf_ram.memory\[112\]\[4\] u_cpu.rf_ram.memory\[113\]\[4\] u_cpu.rf_ram.memory\[114\]\[4\]
+ u_cpu.rf_ram.memory\[115\]\[4\] _01619_ _01620_ _02007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08307_ u_arbiter.i_wb_cpu_rdt\[26\] u_arbiter.i_wb_cpu_rdt\[10\] _01436_ _03888_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09287_ _04484_ _04516_ _04524_ _01246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08453__A2 _04016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06499_ _02790_ _02791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08238_ _03825_ _03826_ _03829_ _03801_ _03832_ _03833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_119_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05929__C _01386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08169_ _03767_ _03768_ _03769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09402__A1 _04468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10200_ _00646_ io_in[4] u_cpu.rf_ram.memory\[127\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07264__I0 _02596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07964__A1 _03551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06767__A2 _02934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10131_ _00577_ io_in[4] u_cpu.rf_ram.memory\[134\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10062_ _00508_ io_in[4] u_cpu.rf_ram.memory\[70\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06519__A2 _02801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07192__A2 _03176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10964_ _10964_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__09602__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10895_ _01324_ io_in[4] u_cpu.rf_ram.memory\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08692__A2 _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06067__I _02516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[66\] u_scanchain_local.module_data_in\[65\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[28\] u_scanchain_local.clk u_scanchain_local.module_data_in\[66\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__09752__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06758__A2 _02934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10329_ _00762_ io_in[4] u_cpu.rf_ram.memory\[117\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05430__A2 _01918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07707__A1 _03357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08755__I0 _02587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05870_ _02309_ _02325_ _01369_ _02352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08380__A1 u_cpu.cpu.immdec.imm30_25\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07183__A2 _03176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05813__S0 _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05194__A1 _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06930__A2 _03031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07540_ _03355_ _03372_ _03378_ _00644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05590__B _01626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06178__S _02578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07471_ _02584_ u_cpu.rf_ram.memory\[12\]\[2\] _03334_ _03337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06422_ _02512_ _02729_ _02736_ _00168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09210_ _04480_ _04470_ _04481_ _01212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06906__S _03021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09141_ u_cpu.rf_ram.memory\[83\]\[1\] _04439_ _04441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06353_ u_cpu.rf_ram.memory\[41\]\[0\] _02697_ _02698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08435__A2 _03776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08406__B _03975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05249__A2 _01739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05304_ _01562_ _01793_ _01582_ _01794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09072_ _04286_ _04399_ _04402_ _01153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06284_ _02502_ _02651_ _02656_ _00110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05749__C _01426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08023_ _03661_ _00845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__06997__A2 _03071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05235_ u_cpu.rf_ram.memory\[36\]\[1\] u_cpu.rf_ram.memory\[37\]\[1\] u_cpu.rf_ram.memory\[38\]\[1\]
+ u_cpu.rf_ram.memory\[39\]\[1\] _01619_ _01620_ _01726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_115_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05166_ u_cpu.rf_ram.memory\[92\]\[0\] u_cpu.rf_ram.memory\[93\]\[0\] u_cpu.rf_ram.memory\[94\]\[0\]
+ u_cpu.rf_ram.memory\[95\]\[0\] _01610_ _01611_ _01658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_115_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07946__A1 _03551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06749__A2 _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09974_ _00428_ io_in[4] u_cpu.rf_ram.memory\[52\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05097_ _01397_ _01589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_58_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08925_ _04321_ _04322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08856_ _03555_ _04271_ _04279_ _01060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08568__S _02445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05056__I _01547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09625__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07174__A2 _03159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08371__A1 _03876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07807_ u_cpu.rf_ram.memory\[117\]\[2\] _03530_ _03533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05804__S0 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08787_ _03543_ _04227_ _04229_ _01041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05999_ _01386_ _01394_ u_cpu.rf_ram_if.genblk1.wtrig0_r _02456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04932__A1 _01434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07738_ _02355_ _02356_ _01369_ _01370_ _03493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__10602__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07669_ u_cpu.rf_ram.memory\[36\]\[7\] _03442_ _03450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08674__A2 _04155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09775__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09408_ _04476_ _04595_ _04599_ _01292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10680_ _01109_ io_in[4] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10752__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09339_ _04482_ _04546_ _04553_ _01269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[4\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06988__A2 _03061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04999__A1 _01445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05660__A2 _02145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10114_ _00560_ io_in[4] u_cpu.rf_ram.memory\[136\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11094_ _11094_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__10132__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10045_ _00491_ io_in[4] u_cpu.rf_ram.memory\[73\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08362__A1 _03876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07165__A2 _03159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10282__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10947_ u_cpu.rf_ram_if.wdata1_r\[1\] io_in[4] u_cpu.rf_ram_if.wdata1_r\[0\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06676__A1 _02750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10878_ _01307_ io_in[4] u_cpu.rf_ram.memory\[25\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08417__A2 _03742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09090__A2 _04409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06979__A2 _03061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05020_ u_arbiter.i_wb_cpu_dbus_adr\[25\] _01457_ _01519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07928__A1 _03551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09648__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05403__A2 _01891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06600__A1 _02746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06971_ _02965_ _03051_ _03057_ _00396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08710_ u_cpu.cpu.ctrl.o_ibus_adr\[25\] _04173_ _04175_ u_cpu.cpu.ctrl.o_ibus_adr\[26\]
+ _04185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_67_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05922_ u_cpu.cpu.ctrl.pc_plus_offset_cy_r _02402_ _02403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__10625__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09690_ _00144_ io_in[4] u_cpu.rf_ram.memory\[41\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08353__A1 _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07156__A2 _03159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05167__A1 _01398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05853_ _01379_ _01382_ _02336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08641_ _03543_ _04145_ _04147_ _00977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09798__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06903__A2 _03012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05784_ _01541_ _02268_ _02269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08572_ u_arbiter.i_wb_cpu_dbus_adr\[7\] u_arbiter.i_wb_cpu_dbus_adr\[6\] _02445_
+ _04108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07523_ u_cpu.rf_ram.memory\[128\]\[6\] _03362_ _03369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10775__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07454_ u_cpu.rf_ram.memory\[130\]\[2\] _03325_ _03328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06405_ _02517_ _02718_ _02726_ _00161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07385_ _03165_ _03285_ _03289_ _00578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08408__A2 u_arbiter.i_wb_cpu_rdt\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10005__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09124_ _04284_ _04429_ _04431_ _01176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07467__I0 _02573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06336_ u_cpu.rf_ram.memory\[51\]\[1\] _02686_ _02688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09081__A2 _04399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09055_ u_cpu.rf_ram.memory\[99\]\[3\] _04389_ _04393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06267_ u_cpu.rf_ram.memory\[42\]\[5\] _02641_ _02647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07467__S _03334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08006_ u_cpu.cpu.bufreg.lsb\[1\] u_cpu.cpu.mem_bytecnt\[1\] _03646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05218_ _01570_ _01708_ _01709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05642__A2 _02128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06198_ _02605_ _00075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10155__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08967__I0 u_arbiter.i_wb_cpu_rdt\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05149_ _01633_ _01635_ _01638_ _01640_ _01628_ _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_116_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09957_ _00411_ io_in[4] u_cpu.rf_ram.memory\[54\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08908_ _04286_ _04309_ _04312_ _01079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09888_ _00342_ io_in[4] u_cpu.rf_ram.memory\[62\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08839_ _02539_ _04197_ _04270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08895__A2 _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05253__S1 _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10801_ _01230_ io_in[4] u_cpu.rf_ram.memory\[10\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08647__A2 _04145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06658__A1 _02750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10732_ _01161_ io_in[4] u_cpu.rf_ram.memory\[105\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10663_ _01092_ io_in[4] u_cpu.rf_ram.memory\[28\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05881__A2 _02313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10594_ _00021_ io_in[4] u_cpu.cpu.alu.add_cy_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08761__S _04208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09072__A2 _04399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06830__A1 _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10648__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[29\] u_arbiter.i_wb_cpu_rdt\[26\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[23\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__07176__I _02516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07386__A2 _03285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09940__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11077_ _11077_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05492__S1 _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08335__A1 _03796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10028_ _00474_ io_in[4] u_cpu.rf_ram.memory\[13\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10798__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06197__I0 _02581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08886__A2 _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05244__S1 _01616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10028__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08638__A2 _04145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06456__S _02756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07310__A2 _03245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07170_ _02506_ _03169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09063__A2 _04389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10178__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06121_ u_cpu.rf_ram.memory\[18\]\[1\] _02551_ _02553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08810__A2 _04242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06052_ _02478_ u_cpu.rf_ram_if.wdata1_r\[5\] _02504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_114_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05003_ _01445_ _01504_ _01505_ u_arbiter.o_wb_cpu_adr\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09811_ _00265_ io_in[4] u_cpu.rf_ram.memory\[75\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09742_ _00196_ io_in[4] u_cpu.rf_ram.memory\[16\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06954_ u_cpu.rf_ram.memory\[57\]\[6\] _03041_ _03048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05483__S1 _01580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07129__A2 _03139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05905_ _02385_ _02386_ _02387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09673_ _00127_ io_in[4] u_cpu.rf_ram.memory\[44\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06885_ u_cpu.rf_ram.memory\[60\]\[7\] _03002_ _03010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05235__S1 _01620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08624_ u_cpu.cpu.bufreg.i_sh_signed _02448_ _02445_ _04135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_54_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05836_ u_cpu.rf_ram_if.rtrig1 _02320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_54_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05767_ _02245_ _02247_ _02249_ _02251_ _01628_ _02252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_78_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08555_ _03549_ _04094_ _04099_ _00939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08629__A2 _02773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07506_ _02516_ _03359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05698_ _01614_ _02183_ _01654_ _02184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08486_ u_cpu.cpu.immdec.imm19_12_20\[5\] _04016_ _04049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07301__A2 _03235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07437_ _03163_ _03315_ _03318_ _00601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05863__A2 _02338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09054__A2 _04389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09813__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07368_ u_cpu.rf_ram.memory\[135\]\[4\] _03275_ _03280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09107_ u_cpu.rf_ram.memory\[106\]\[2\] _04419_ _04422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07065__A1 _02577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06319_ u_cpu.rf_ram.memory\[44\]\[3\] _02673_ _02677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07299_ _03169_ _03235_ _03241_ _00540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09038_ _04288_ _04379_ _04383_ _01138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09963__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07368__A2 _03275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11000_ _11000_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_105_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05379__A1 _01406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05918__A3 _02372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10940__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05474__S1 _01557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08317__A1 _03831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05226__S1 _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07540__A2 _03372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09293__A2 _04526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10320__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10715_ _01144_ io_in[4] u_cpu.rf_ram.memory\[99\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10646_ _01075_ io_in[4] u_cpu.rf_ram.memory\[95\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09045__A2 _04379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10577_ _01007_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10470__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05606__A2 _02092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06803__I _02501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08223__C _03810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08308__A1 _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05582__C _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05790__A1 _01398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05217__S1 _01574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06670_ _02744_ _02884_ _02887_ _00265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05154__I _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07531__A2 _03372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05621_ _02101_ _02103_ _02105_ _02107_ _01426_ _02108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_24_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05393__I1 u_cpu.rf_ram.memory\[29\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08340_ _02768_ _03914_ _03919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05552_ _01684_ _02039_ _01418_ _02040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06186__S _02578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09836__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09284__A2 _04516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07295__A1 _03165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08271_ _03767_ _03861_ _03862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05483_ u_cpu.rf_ram.memory\[24\]\[4\] u_cpu.rf_ram.memory\[25\]\[4\] u_cpu.rf_ram.memory\[26\]\[4\]
+ u_cpu.rf_ram.memory\[27\]\[4\] _01578_ _01580_ _01971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_20_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07222_ _03163_ _03196_ _03199_ _00505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10813__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09036__A2 _04379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06914__S _03021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07047__A1 _02969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07153_ _02481_ _03157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09986__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07598__A2 _03402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08795__A1 _03551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06104_ _02487_ _02541_ _02543_ _00043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08414__B _03983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07084_ u_cpu.rf_ram.memory\[142\]\[0\] _03119_ _03120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06035_ _02460_ u_cpu.rf_ram_if.wdata0_r\[2\] _02489_ _02490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06270__A2 _02641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08547__A1 _03539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05773__B _01416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06022__A2 _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07986_ _03555_ _03626_ _03634_ _00835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07770__A2 _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09725_ _00179_ io_in[4] u_cpu.rf_ram.memory\[4\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06937_ _02967_ _03031_ _03038_ _00381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05208__S1 _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09656_ _00110_ io_in[4] u_cpu.rf_ram.memory\[46\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08576__S _02445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06868_ _02969_ _02992_ _03000_ _00350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05064__I _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07522__A2 _03362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10343__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08607_ u_arbiter.i_wb_cpu_dbus_adr\[24\] u_arbiter.i_wb_cpu_dbus_adr\[23\] _04115_
+ _04126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_63_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05819_ _01406_ _02254_ _02303_ _00007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_70_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09587_ _00041_ io_in[4] u_cpu.rf_ram.memory\[21\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06799_ _02959_ _02955_ _02960_ _00321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08538_ u_cpu.rf_ram.memory\[32\]\[5\] _04084_ _04090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09275__A2 _04516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06089__A2 _02530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07286__A1 _02602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08469_ _04029_ _04004_ _04032_ _03782_ _04033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10493__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10500_ _00933_ io_in[4] u_cpu.rf_ram.memory\[32\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09027__A2 _04369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10431_ _00864_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07589__A2 _03402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10362_ _00795_ io_in[4] u_cpu.rf_ram.memory\[8\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06261__A2 _02641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05695__S1 _01620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10293_ _00726_ io_in[4] u_cpu.rf_ram.memory\[90\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[3\]_D u_arbiter.i_wb_cpu_rdt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09709__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07210__A1 _03169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07761__A2 _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09859__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07513__A2 _03362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05524__A1 _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10836__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09266__A2 _04506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07277__A1 _03165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09018__A2 _04369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07029__A1 _02969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10629_ _01058_ io_in[4] u_cpu.rf_ram.memory\[97\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10216__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05686__S1 _01549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08529__A1 _03539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06004__A2 _02460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07840_ u_cpu.rf_ram.memory\[120\]\[6\] _03541_ _03554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07752__A2 _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10366__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07771_ u_cpu.rf_ram.memory\[35\]\[2\] _03510_ _03513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04983_ u_cpu.cpu.ctrl.o_ibus_adr\[16\] _01488_ _01491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_49_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09510_ u_cpu.rf_ram.memory\[100\]\[1\] _04654_ _04656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06722_ _02742_ _02914_ _02916_ _00288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07504__A2 _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09441_ u_cpu.rf_ram.memory\[25\]\[2\] _04615_ _04618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06653_ u_cpu.rf_ram.memory\[76\]\[3\] _02874_ _02878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05604_ _01589_ _02090_ _02091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09372_ _04575_ _01280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09257__A2 _04506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06584_ _02748_ _02834_ _02839_ _00227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08323_ _03897_ _03903_ _03904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07268__A1 _02638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05535_ _01667_ _02022_ _02023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05818__A2 _02302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08254_ u_arbiter.i_wb_cpu_rdt\[20\] u_arbiter.i_wb_cpu_rdt\[4\] _01437_ _03846_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05466_ _01945_ _01954_ _01955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09009__A2 _04359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07205_ u_cpu.rf_ram.memory\[71\]\[3\] _03186_ _03190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08185_ _02765_ u_arbiter.i_wb_cpu_rdt\[13\] _03784_ _03785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05397_ _01879_ _01881_ _01883_ _01885_ _01426_ _01886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_07136_ _02577_ _02660_ _03148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06243__A2 _02628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07067_ _03110_ _00439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05677__S1 _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06018_ _02474_ _02475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07475__S _03334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07991__A2 _03636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10709__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05429__S1 _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07743__A2 _02395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07969_ _02561_ _02821_ _03625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09708_ _00162_ io_in[4] u_cpu.rf_ram.memory\[47\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10980_ _10980_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__10859__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09496__A2 _04644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09639_ _00093_ io_in[4] u_cpu.rf_ram.memory\[78\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05678__B _01626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10239__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05690__B1 _02173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10414_ _00847_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05397__C _01426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09420__A2 _04605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06234__A2 _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10345_ _00778_ io_in[4] u_cpu.rf_ram.memory\[118\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05668__S1 _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07982__A2 _03626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10389__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10276_ _00709_ io_in[4] u_cpu.cpu.state.o_cnt_r\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09184__A1 _04290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[11\] u_arbiter.i_wb_cpu_rdt\[8\] io_in[3] u_arbiter.i_wb_cpu_dbus_dat\[5\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__08501__C _03791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09681__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08931__A1 _04286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07498__A1 u_cpu.rf_ram.memory\[22\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08998__A1 _04284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05320_ _01609_ _01809_ _01810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06464__S _02756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08462__A3 _03768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05251_ u_cpu.rf_ram.memory\[124\]\[1\] u_cpu.rf_ram.memory\[125\]\[1\] u_cpu.rf_ram.memory\[126\]\[1\]
+ u_cpu.rf_ram.memory\[127\]\[1\] _01545_ _01642_ _01742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07670__A1 _03359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06473__A2 _02769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05182_ _01667_ _01673_ _01674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09411__A2 _04595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06225__A2 _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05659__S1 _01580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09990_ _00444_ io_in[4] u_cpu.rf_ram.memory\[15\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07973__A2 _03626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08941_ _04296_ _04322_ _04330_ _01094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08872_ u_cpu.rf_ram.memory\[94\]\[4\] _04282_ _04291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07725__A2 _03475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08922__A1 _01437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07823_ _03539_ _03541_ _03542_ _00764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07754_ _03349_ _03500_ _03503_ _00734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_04966_ u_cpu.cpu.ctrl.o_ibus_adr\[12\] _01476_ _01478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_93_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07489__A1 u_cpu.rf_ram.memory\[22\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06705_ u_cpu.rf_ram.memory\[68\]\[2\] _02904_ _02907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08686__B1 _04157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07685_ u_cpu.rf_ram_if.rgnt _03460_ _02433_ _01429_ _03461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_52_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04897_ u_cpu.cpu.immdec.imm19_12_20\[6\] _01368_ _01423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09424_ _04474_ _04605_ _04608_ _01299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06636_ _02746_ _02864_ _02868_ _00250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_u_scanchain_local.scan_flop\[27\]_D u_arbiter.i_wb_cpu_rdt\[24\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06161__A1 _02539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09355_ _04480_ _04556_ _04562_ _01276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06567_ _02750_ _02823_ _02829_ _00220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08306_ _03555_ _03879_ _03887_ _00902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05518_ _01645_ _02005_ _01648_ _02006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_139_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09286_ u_cpu.rf_ram.memory\[110\]\[7\] _04516_ _04524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06498_ _02528_ _02612_ _02790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05498__B _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08237_ _03782_ _03804_ _03831_ _03832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05449_ _01553_ _01937_ _01565_ _01938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_101_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08168_ u_arbiter.i_wb_cpu_rdt\[15\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\]
+ _01436_ _03768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09402__A2 _04595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10531__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06216__A2 _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07119_ _03138_ _03139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08099_ u_arbiter.i_wb_cpu_rdt\[24\] _03669_ _03715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07964__A2 _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10130_ _00576_ io_in[4] u_cpu.rf_ram.memory\[134\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05975__A1 u_cpu.cpu.decode.opcode\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09166__A1 _04290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10061_ _00507_ io_in[4] u_cpu.rf_ram.memory\[70\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10681__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07716__A2 _03475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09469__A2 _04625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10963_ _10963_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__04950__A2 _01457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[18\]_D u_arbiter.i_wb_cpu_rdt\[15\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06152__A1 _02512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10894_ _01323_ io_in[4] u_cpu.rf_ram.memory\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10061__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07652__A1 _03359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[59\] u_scanchain_local.module_data_in\[58\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[21\] u_scanchain_local.clk u_scanchain_local.module_data_in\[59\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_138_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07955__A2 _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10328_ _00761_ io_in[4] u_cpu.rf_ram.memory\[117\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05510__S0 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10259_ _00692_ io_in[4] u_cpu.rf_ram.memory\[37\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07707__A2 _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[32\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08904__A1 _04280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05569__I1 u_cpu.rf_ram.memory\[29\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05813__S1 _01574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06391__A1 _02482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08668__B1 _04157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[10\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08132__A2 _03731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10404__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07470_ _03336_ _00616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05162__I _01564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06421_ u_cpu.rf_ram.memory\[47\]\[6\] _02729_ _02736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09577__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09140_ _04280_ _04439_ _04440_ _01183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06352_ _02696_ _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_u_scanchain_local.scan_flop\[25\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10554__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05303_ u_cpu.rf_ram.memory\[16\]\[2\] u_cpu.rf_ram.memory\[17\]\[2\] u_cpu.rf_ram.memory\[18\]\[2\]
+ u_cpu.rf_ram.memory\[19\]\[2\] _01578_ _01580_ _01793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_06283_ u_cpu.rf_ram.memory\[46\]\[4\] _02651_ _02656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06446__A2 _02740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09071_ u_cpu.rf_ram.memory\[79\]\[2\] _04399_ _04402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08022_ u_arbiter.i_wb_cpu_rdt\[1\] _02781_ _03660_ _03661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05234_ _01614_ _01724_ _01605_ _01725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09396__A1 _03812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05165_ _01422_ _01641_ _01656_ _01657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_116_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07946__A2 _03606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09973_ _00427_ io_in[4] u_cpu.rf_ram.memory\[52\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05096_ _01576_ _01583_ _01585_ _01587_ _01426_ _01588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__05501__S0 _01623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05957__A1 _01403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09148__A1 _04290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08924_ _02528_ _02671_ _04321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08855_ u_cpu.rf_ram.memory\[97\]\[7\] _04271_ _04279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07806_ _03347_ _03530_ _03532_ _00757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05804__S1 _01549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08786_ u_cpu.rf_ram.memory\[93\]\[1\] _04227_ _04229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05185__A2 _01672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05998_ _02431_ _02455_ _02332_ u_arbiter.i_wb_cpu_dbus_sel\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07737_ _01408_ _02332_ _03488_ _03490_ _03492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_44_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04949_ _01463_ _01464_ _01465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10084__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07668_ _03357_ _03442_ _03449_ _00701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08584__S _02445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06134__A1 _02517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09407_ u_cpu.rf_ram.memory\[27\]\[3\] _04595_ _04599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06619_ u_cpu.rf_ram.memory\[77\]\[4\] _02854_ _02859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07599_ _02706_ _02821_ _03411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09338_ u_cpu.rf_ram.memory\[87\]\[6\] _04546_ _04553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07634__A1 _03359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06437__A2 _02740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09269_ _04484_ _04506_ _04514_ _01238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09387__A1 _02339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[55\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07937__A2 _03606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05948__A1 _02320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10113_ _00559_ io_in[4] u_cpu.rf_ram.memory\[136\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11093_ _11093_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_1_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08759__S _04208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10044_ _00490_ io_in[4] u_cpu.rf_ram.memory\[73\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_scanchain_local.scan_flop\[4\] u_arbiter.i_wb_cpu_rdt\[1\] io_in[3] u_arbiter.i_wb_cpu_dbus_sel\[2\]
+ u_scanchain_local.clk u_arbiter.i_wb_cpu_rdt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_75_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10427__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06373__A1 _02482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09311__A1 _04472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10946_ _01365_ io_in[4] u_cpu.rf_ram_if.rcnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10577__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06676__A2 _02884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10877_ _01306_ io_in[4] u_cpu.rf_ram.memory\[25\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06920__I0 _02599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06806__I _02506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06428__A2 _02740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07928__A2 _03596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05939__A1 _02320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06600__A2 _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06970_ u_cpu.rf_ram.memory\[56\]\[5\] _03051_ _03057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05921_ u_arbiter.i_wb_cpu_ibus_adr\[0\] _02401_ _02402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08353__A2 _03926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08640_ u_cpu.rf_ram.memory\[30\]\[1\] _04145_ _04147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05852_ _01370_ _02331_ _02333_ _02335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06364__A1 _02507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05798__S0 _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08571_ _04107_ _00947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_81_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05783_ u_cpu.rf_ram.memory\[112\]\[7\] u_cpu.rf_ram.memory\[113\]\[7\] u_cpu.rf_ram.memory\[114\]\[7\]
+ u_cpu.rf_ram.memory\[115\]\[7\] _01619_ _01620_ _02268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_35_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08105__A2 _03718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07522_ _03355_ _03362_ _03368_ _00636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06116__A1 _02517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07453_ _03161_ _03325_ _03327_ _00608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06667__A2 _02884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06404_ u_cpu.rf_ram.memory\[48\]\[7\] _02718_ _02726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07384_ u_cpu.rf_ram.memory\[134\]\[3\] _03285_ _03289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09123_ u_cpu.rf_ram.memory\[107\]\[1\] _04429_ _04431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07616__A1 _03359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06419__A2 _02729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06335_ _02482_ _02686_ _02687_ _00130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09054_ _04286_ _04389_ _04392_ _01145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06266_ _02502_ _02641_ _02646_ _00102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07092__A2 _03119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08005_ u_cpu.cpu.bufreg.lsb\[1\] u_cpu.cpu.mem_bytecnt\[1\] u_cpu.cpu.mem_bytecnt\[0\]
+ u_cpu.cpu.bufreg.lsb\[0\] _03645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__09369__A1 _01375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09369__B2 _01385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05217_ u_cpu.rf_ram.memory\[28\]\[1\] u_cpu.rf_ram.memory\[29\]\[1\] u_cpu.rf_ram.memory\[30\]\[1\]
+ u_cpu.rf_ram.memory\[31\]\[1\] _01572_ _01574_ _01708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_06197_ _02581_ u_cpu.rf_ram.memory\[7\]\[1\] _02603_ _02605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07919__A2 _03596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04850__A1 _01373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08041__A1 u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05148_ _01601_ _01639_ _01626_ _01640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09956_ _00410_ io_in[4] u_cpu.rf_ram.memory\[54\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05079_ _01544_ _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_131_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08329__C1 _03826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08907_ u_cpu.rf_ram.memory\[96\]\[2\] _04309_ _04312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09887_ _00341_ io_in[4] u_cpu.rf_ram.memory\[62\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09742__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09541__A1 _04484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08344__A2 _03914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08838_ _02525_ _04237_ _04268_ _04269_ _01052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_45_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05789__S0 _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08769_ _04219_ _01033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10800_ _01229_ io_in[4] u_cpu.rf_ram.memory\[10\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09892__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10731_ _01160_ io_in[4] u_cpu.rf_ram.memory\[105\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06658__A2 _02874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10662_ _01091_ io_in[4] u_cpu.rf_ram.memory\[28\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10593_ _01023_ io_in[4] u_cpu.rf_ram.memory\[109\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08280__A1 _03791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06830__A2 _02972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06594__A1 _02738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05397__A2 _01881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11076_ _11076_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_62_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08335__A2 _03914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10027_ _00473_ io_in[4] u_cpu.rf_ram.memory\[13\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06897__A2 _03012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08099__A1 u_arbiter.i_wb_cpu_rdt\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10929_ _01357_ io_in[4] u_cpu.rf_ram.memory\[23\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06649__A2 _02874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08237__B _03831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06120_ _02482_ _02551_ _02552_ _00050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08271__A1 _03767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09615__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06051_ _02477_ _02502_ _02503_ _00030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06821__A2 _02972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05002_ u_arbiter.i_wb_cpu_dbus_adr\[21\] _01457_ _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09765__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09810_ _00264_ io_in[4] u_cpu.rf_ram.memory\[75\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09741_ _00195_ io_in[4] u_cpu.rf_ram.memory\[16\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06953_ _02965_ _03041_ _03047_ _00388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10742__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09523__A1 _04484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05904_ u_arbiter.i_wb_cpu_dbus_dat\[0\] u_arbiter.i_wb_cpu_dbus_dat\[8\] u_arbiter.i_wb_cpu_dbus_dat\[16\]
+ u_arbiter.i_wb_cpu_dbus_dat\[24\] u_cpu.cpu.bufreg.lsb\[0\] u_cpu.cpu.bufreg.lsb\[1\]
+ _02386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA_u_scanchain_local.scan_flop\[3\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09672_ _00126_ io_in[4] u_cpu.rf_ram.memory\[44\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08198__I _03796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06884_ _02967_ _03002_ _03009_ _00357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06337__A1 _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06188__I1 u_cpu.cpu.o_wdata0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08623_ _04133_ _02445_ _04134_ _00972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05835_ _02311_ _02315_ _02316_ _02318_ _02319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08554_ u_cpu.rf_ram.memory\[31\]\[4\] _04094_ _04099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05766_ _01645_ _02250_ _01626_ _02251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07137__I0 _02573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10892__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07830__I _02496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07505_ _03357_ _03345_ _03358_ _00629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07837__A1 u_cpu.rf_ram.memory\[120\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08485_ u_cpu.cpu.immdec.imm19_12_20\[6\] _02768_ _04048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05697_ u_cpu.rf_ram.memory\[116\]\[6\] u_cpu.rf_ram.memory\[117\]\[6\] u_cpu.rf_ram.memory\[118\]\[6\]
+ u_cpu.rf_ram.memory\[119\]\[6\] _01623_ _01624_ _02183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07436_ u_cpu.rf_ram.memory\[131\]\[2\] _03315_ _03318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10122__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07367_ _03165_ _03275_ _03279_ _00570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09106_ _04284_ _04419_ _04421_ _01168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06318_ _02492_ _02673_ _02676_ _00124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07065__A2 _02727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07298_ u_cpu.rf_ram.memory\[39\]\[5\] _03235_ _03241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09037_ u_cpu.rf_ram.memory\[104\]\[3\] _04379_ _04383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06249_ _02512_ _02628_ _02635_ _00096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10272__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08014__A1 _03653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05379__A2 _01819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06576__A1 _02738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09939_ _00393_ io_in[4] u_cpu.rf_ram.memory\[56\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08317__A2 _03776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06328__A1 _02517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06879__A2 _03002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10714_ _01143_ io_in[4] u_cpu.rf_ram.memory\[99\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08772__S _04217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09638__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10645_ _01074_ io_in[4] u_cpu.rf_ram.memory\[95\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10615__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08253__A1 _01408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10576_ _01006_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05067__A1 _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09788__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[41\] u_scanchain_local.module_data_in\[40\] io_in[3]
+ u_arbiter.o_wb_cpu_adr\[3\] u_scanchain_local.clk u_scanchain_local.module_data_in\[41\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_127_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08005__A1 u_cpu.cpu.bufreg.lsb\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10765__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08556__A2 _04094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06567__A1 _02750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09505__A1 _04484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11059_ _11059_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_77_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08947__S _04331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05620_ _01614_ _02106_ _01654_ _02107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_58_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05542__A2 _02025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10145__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05551_ u_cpu.rf_ram.memory\[132\]\[4\] u_cpu.rf_ram.memory\[133\]\[4\] u_cpu.rf_ram.memory\[134\]\[4\]
+ u_cpu.rf_ram.memory\[135\]\[4\] _01687_ _01688_ _02039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_60_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08270_ _03768_ _03802_ _03861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07295__A2 _03235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08492__A1 _04024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05482_ _01570_ _01969_ _01970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07221_ u_cpu.rf_ram.memory\[70\]\[2\] _03196_ _03199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10295__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08244__A1 _03761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07152_ _03156_ _00478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07047__A2 _03091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06103_ u_cpu.rf_ram.memory\[81\]\[1\] _02541_ _02543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08795__A2 _04227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07083_ _03118_ _03119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06034_ _02478_ u_cpu.rf_ram_if.wdata1_r\[2\] _02489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_133_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08547__A2 _04094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06558__A1 u_cpu.rf_ram.memory\[119\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05605__I0 u_cpu.rf_ram.memory\[120\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07985_ u_cpu.rf_ram.memory\[116\]\[7\] _03626_ _03634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09724_ _00178_ io_in[4] u_cpu.rf_ram.memory\[4\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06936_ u_cpu.rf_ram.memory\[58\]\[6\] _03031_ _03038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09655_ _00109_ io_in[4] u_cpu.rf_ram.memory\[46\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06867_ u_cpu.rf_ram.memory\[61\]\[7\] _02992_ _03000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08606_ _04125_ _00964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05818_ _02293_ _02302_ _02303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09586_ _00040_ io_in[4] u_cpu.rf_ram.memory\[21\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06798_ u_cpu.rf_ram.memory\[29\]\[2\] _02955_ _02960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06730__A1 _02750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08537_ _03549_ _04084_ _04089_ _00931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05749_ _02227_ _02229_ _02231_ _02233_ _01426_ _02234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__10638__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08468_ _03999_ _03988_ _04030_ _04031_ _03801_ _04032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__07286__A2 _02639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05080__I _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05297__A1 _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07419_ _03163_ _03305_ _03308_ _00593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08399_ _03969_ _03970_ _03906_ _03971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_13_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09930__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10430_ _00863_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07038__A2 _03091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10788__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08786__A2 _04227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10361_ _00794_ io_in[4] u_cpu.rf_ram.memory\[8\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10292_ _00725_ io_in[4] u_cpu.rf_ram.memory\[90\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08538__A2 _04084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10018__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07210__A2 _03186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10168__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08710__A2 _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05524__A2 _02002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07277__A2 _03225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05288__A1 _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10628_ _01057_ io_in[4] u_cpu.rf_ram.memory\[97\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08226__A1 _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07029__A2 _03081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10559_ _00989_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06788__A1 _02754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08529__A2 _04084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05460__A1 _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07201__A2 _03186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07770_ _03347_ _03510_ _03512_ _00741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_04982_ u_cpu.cpu.ctrl.o_ibus_adr\[16\] _01488_ _01490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09803__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06721_ u_cpu.rf_ram.memory\[67\]\[1\] _02914_ _02916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09440_ _04472_ _04615_ _04617_ _01306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_64_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06652_ _02744_ _02874_ _02877_ _00257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06197__S _02603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06712__A1 _02750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05603_ u_cpu.rf_ram.memory\[124\]\[5\] u_cpu.rf_ram.memory\[125\]\[5\] u_cpu.rf_ram.memory\[126\]\[5\]
+ u_cpu.rf_ram.memory\[127\]\[5\] _01545_ _01642_ _02090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_91_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05071__S0 _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09371_ _04574_ u_cpu.cpu.genblk3.csr.mcause3_0\[1\] _04568_ _04575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_52_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06583_ u_cpu.rf_ram.memory\[129\]\[4\] _02834_ _02839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09953__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08322_ _03861_ _03899_ _03902_ _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_21_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05114__B _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05534_ u_cpu.rf_ram.memory\[64\]\[4\] u_cpu.rf_ram.memory\[65\]\[4\] u_cpu.rf_ram.memory\[66\]\[4\]
+ u_cpu.rf_ram.memory\[67\]\[4\] _01571_ _01668_ _02022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08465__A1 _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07268__A2 _02832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05279__A1 _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08253_ _01408_ _03740_ _03845_ _00891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10930__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05465_ _01947_ _01949_ _01951_ _01953_ _01404_ _01954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_119_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07204_ _03163_ _03186_ _03189_ _00497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08217__A1 _03796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08184_ _01435_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[13\] _03784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05396_ _01542_ _01884_ _01418_ _01885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_134_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07135_ _02969_ _03139_ _03147_ _00470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07066_ _02573_ u_cpu.rf_ram.memory\[15\]\[0\] _03109_ _03110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07440__A2 _03315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05451__A1 _01667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06017_ u_cpu.cpu.immdec.imm11_7\[3\] _02470_ _02473_ _02474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_82_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10310__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05203__A1 _01406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08940__A2 _04322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07968_ _03555_ _03616_ _03624_ _00827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08587__S _04115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06951__A1 _02963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06919_ _03028_ _00373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09707_ _00161_ io_in[4] u_cpu.rf_ram.memory\[48\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_u_scanchain_local.scan_flop\[6\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07899_ _02573_ u_cpu.rf_ram.memory\[11\]\[0\] _03586_ _03587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10460__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09638_ _00092_ io_in[4] u_cpu.rf_ram.memory\[78\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09569_ u_cpu.rf_ram_if.rcnt\[1\] u_cpu.rf_ram_if.rcnt\[0\] _04688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_31_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08456__B2 _03840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08208__A1 _03798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10413_ _00846_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10344_ _00777_ io_in[4] u_cpu.rf_ram.memory\[118\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05442__A1 _01609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05694__B _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10275_ _00708_ io_in[4] u_cpu.cpu.state.o_cnt_r\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09826__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09184__A2 _04459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08931__A2 _04322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10803__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09976__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07498__A2 _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06809__I _02511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10953__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08447__A1 _02305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08998__A2 _04359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05250_ _01734_ _01736_ _01738_ _01740_ _01628_ _01741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_31_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07670__A2 _03442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05681__A1 _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05181_ u_cpu.rf_ram.memory\[72\]\[0\] u_cpu.rf_ram.memory\[73\]\[0\] u_cpu.rf_ram.memory\[74\]\[0\]
+ u_cpu.rf_ram.memory\[75\]\[0\] _01571_ _01668_ _01673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_128_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08080__C1 _03676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07422__A2 _03305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10333__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08940_ u_cpu.rf_ram.memory\[28\]\[7\] _04322_ _04330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09175__A2 _04459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08871_ _02501_ _04290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_111_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07186__A1 _03163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07822_ u_cpu.rf_ram.memory\[120\]\[0\] _03541_ _03542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10483__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06933__A1 _02963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05292__S0 _01546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07753_ u_cpu.rf_ram.memory\[92\]\[2\] _03500_ _03503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04965_ _01443_ _01474_ _01476_ _01477_ u_arbiter.o_wb_cpu_adr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_38_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06704_ _02742_ _02904_ _02906_ _00280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_93_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07489__A2 _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08686__A1 u_cpu.cpu.ctrl.o_ibus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07684_ _02783_ _03460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08686__B2 u_cpu.cpu.ctrl.o_ibus_adr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04896_ _01421_ _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_92_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09423_ u_cpu.rf_ram.memory\[26\]\[2\] _04605_ _04608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06635_ u_cpu.rf_ram.memory\[74\]\[3\] _02864_ _02868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06161__A2 _02577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09354_ u_cpu.rf_ram.memory\[88\]\[5\] _04556_ _04562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06566_ u_cpu.rf_ram.memory\[119\]\[5\] _02823_ _02829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08438__A1 _03754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09486__I0 _02599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08305_ u_cpu.rf_ram.memory\[114\]\[7\] _03879_ _03887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05517_ u_cpu.rf_ram.memory\[120\]\[4\] u_cpu.rf_ram.memory\[121\]\[4\] u_cpu.rf_ram.memory\[122\]\[4\]
+ u_cpu.rf_ram.memory\[123\]\[4\] _01646_ _01603_ _02005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08989__A2 _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09285_ _04482_ _04516_ _04523_ _01245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06497_ _02784_ _02789_ _00190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08236_ _03830_ _03831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05448_ u_cpu.rf_ram.memory\[68\]\[3\] u_cpu.rf_ram.memory\[69\]\[3\] u_cpu.rf_ram.memory\[70\]\[3\]
+ u_cpu.rf_ram.memory\[71\]\[3\] _01555_ _01652_ _01937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09238__I0 _02581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07661__A2 _03442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05672__A1 _01609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08167_ _02765_ u_arbiter.i_wb_cpu_rdt\[14\] _03766_ _03767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05379_ _01406_ _01819_ _01868_ _00002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_134_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07118_ _02671_ _02832_ _03138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09849__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08098_ _03713_ _03714_ _00867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07049_ _02573_ u_cpu.rf_ram.memory\[9\]\[0\] _03100_ _03101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10826__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05975__A2 _02313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09166__A2 _04449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10060_ _00506_ io_in[4] u_cpu.rf_ram.memory\[70\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09999__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08913__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05283__S0 _01680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10962_ _10962_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_29_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10893_ _01322_ io_in[4] u_cpu.rf_ram.memory\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06152__A2 _02563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10206__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08429__A1 _01436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05689__B _01626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07652__A2 _03432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08780__S _04217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10356__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05663__A1 _01589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05201__C _01404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07404__A2 _03295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10327_ _00760_ io_in[4] u_cpu.rf_ram.memory\[117\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05510__S1 _01549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09157__A2 _04449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10258_ _00691_ io_in[4] u_cpu.rf_ram.memory\[37\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08904__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10189_ _00635_ io_in[4] u_cpu.rf_ram.memory\[128\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05718__A2 _02199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05569__I2 u_cpu.rf_ram.memory\[30\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05274__S0 _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06391__A2 _02718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08955__S _04331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07340__A1 _02810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06143__A2 _02563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06420_ _02507_ _02729_ _02735_ _00167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06351_ _02639_ _02695_ _02696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05302_ _01570_ _01791_ _01792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09070_ _04284_ _04399_ _04401_ _01152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06282_ _02497_ _02651_ _02655_ _00109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07643__A2 _03432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08021_ _03656_ _03658_ _02781_ _03659_ _03660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__05654__A1 _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05233_ u_cpu.rf_ram.memory\[44\]\[1\] u_cpu.rf_ram.memory\[45\]\[1\] u_cpu.rf_ram.memory\[46\]\[1\]
+ u_cpu.rf_ram.memory\[47\]\[1\] _01615_ _01616_ _01724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_128_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10849__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05164_ _01644_ _01649_ _01651_ _01655_ _01607_ _01656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_143_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06454__I0 _02581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09972_ _00426_ io_in[4] u_cpu.rf_ram.memory\[52\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05095_ _01542_ _01586_ _01418_ _01587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_131_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05501__S1 _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09148__A2 _04439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08923_ _01428_ _04320_ _01086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_130_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08854_ _03553_ _04271_ _04278_ _01059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05709__A2 _02190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07833__I _02501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05265__S0 _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07805_ u_cpu.rf_ram.memory\[117\]\[1\] _03530_ _03532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08785_ _03539_ _04227_ _04228_ _01040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05997_ u_cpu.cpu.bufreg.lsb\[0\] _02431_ _02332_ u_arbiter.i_wb_cpu_dbus_sel\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06382__A2 _02708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10229__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07736_ _03488_ _03490_ _03491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_04948_ _01461_ _01462_ _01464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_66_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09320__A2 _04536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07667_ u_cpu.rf_ram.memory\[36\]\[6\] _03442_ _03449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04879_ _01402_ _01404_ _01405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_26_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06134__A2 _02551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07331__A1 _03165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06618_ _02746_ _02854_ _02858_ _00242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09406_ _04474_ _04595_ _04598_ _01291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07598_ _03359_ _03402_ _03410_ _00670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10379__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09337_ _04480_ _04546_ _04552_ _01268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06549_ u_cpu.rf_ram.memory\[40\]\[6\] _02812_ _02819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09671__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09268_ u_cpu.rf_ram.memory\[85\]\[7\] _04506_ _04514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07634__A2 _03422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05645__A1 _01542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08219_ _01372_ _03798_ _03762_ _03816_ _03817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06693__I0 _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09199_ _02491_ _04474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09387__A2 _03454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__04860__C _01385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09139__A2 _04439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10112_ _00558_ io_in[4] u_cpu.rf_ram.memory\[49\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11092_ _11092_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_121_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08347__B1 _03818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10043_ _00489_ io_in[4] u_cpu.rf_ram.memory\[73\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08898__A1 _04294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07570__A1 _03349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06373__A2 _02708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09311__A2 _04536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10945_ u_cpu.rf_ram_if.rtrig0 io_in[4] u_cpu.rf_ram_if.rtrig1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07322__A1 _02539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06125__A2 _02551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07873__A2 _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10876_ _01305_ io_in[4] u_cpu.rf_ram.memory\[25\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05884__A1 _02305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07625__A2 _03422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08822__A1 _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05636__A1 _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09378__A2 _04568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07389__A1 _03169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05495__S0 _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05920_ _01374_ _02306_ _01381_ _01378_ _02400_ _02401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_67_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09550__A2 _04674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05851_ _02332_ _02333_ _02334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06364__A2 _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05798__S1 _01668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08570_ u_arbiter.i_wb_cpu_dbus_adr\[6\] u_arbiter.i_wb_cpu_dbus_adr\[5\] _02445_
+ _04107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05782_ _01601_ _02266_ _01605_ _02267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_19_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07521_ u_cpu.rf_ram.memory\[128\]\[5\] _03362_ _03368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09302__A2 _04526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10521__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06116__A2 _02541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07313__A1 _03165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07452_ u_cpu.rf_ram.memory\[130\]\[1\] _03325_ _03327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09694__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05901__I _02313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05875__A1 _01369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06403_ _02512_ _02718_ _02725_ _00160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08417__C _03818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07383_ _03163_ _03285_ _03288_ _00577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09122_ _04280_ _04429_ _04430_ _01175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10671__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06334_ u_cpu.rf_ram.memory\[51\]\[0\] _02686_ _02687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07616__A2 _03412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05627__A1 _01667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09053_ u_cpu.rf_ram.memory\[99\]\[2\] _04389_ _04392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06265_ u_cpu.rf_ram.memory\[42\]\[4\] _02641_ _02646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08004_ _03555_ _03636_ _03644_ _00843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09369__A2 _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05216_ _01562_ _01706_ _01582_ _01707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06196_ _02604_ _00074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04850__A2 _01375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05147_ u_cpu.rf_ram.memory\[96\]\[0\] u_cpu.rf_ram.memory\[97\]\[0\] u_cpu.rf_ram.memory\[98\]\[0\]
+ u_cpu.rf_ram.memory\[99\]\[0\] _01602_ _01579_ _01639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08041__A2 _02774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06052__A1 _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05486__S0 _01590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09955_ _00409_ io_in[4] u_cpu.rf_ram.memory\[54\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05078_ _01398_ _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_106_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08329__B1 _03769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08329__C2 _03744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08906_ _04284_ _04309_ _04311_ _01078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05792__B _01648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10051__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09886_ _00340_ io_in[4] u_cpu.rf_ram.memory\[62\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09541__A2 _04664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08837_ u_cpu.cpu.immdec.imm30_25\[0\] _03798_ _04237_ _04269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07552__A1 _03349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06355__A2 _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05789__S1 _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08595__S _04115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08768_ _02581_ u_cpu.rf_ram.memory\[2\]\[1\] _04217_ _04219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07719_ _03351_ _03475_ _03479_ _00722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06107__A2 _02541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07304__A1 _02695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08699_ _04179_ _01003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_54_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10730_ _01159_ io_in[4] u_cpu.rf_ram.memory\[105\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07855__A2 _03558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08327__C _03800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05866__A1 _01393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10661_ _01090_ io_in[4] u_cpu.rf_ram.memory\[28\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07607__A2 _03412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10592_ _01022_ io_in[4] u_cpu.rf_ram.memory\[109\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08804__A1 _03860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[22\]_SE io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05618__A1 _01609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05477__S0 _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06594__A2 _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11075_ _11075_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_23_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[24\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10026_ _00472_ io_in[4] u_cpu.rf_ram.memory\[13\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09532__A2 _04664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10544__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06346__A2 _02686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05207__B _01417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[39\]_CLK u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08099__A2 _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10694__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10928_ _01356_ io_in[4] u_cpu.rf_ram.memory\[23\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05857__A1 _02337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10859_ _01288_ io_in[4] u_cpu.cpu.genblk3.csr.o_new_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_75_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06282__A1 _02497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06050_ u_cpu.rf_ram.memory\[82\]\[4\] _02477_ _02503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05001_ u_cpu.cpu.ctrl.o_ibus_adr\[21\] _01503_ _01504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xu_scanchain_local.output_buffers\[3\] u_scanchain_local.clk u_scanchain_local.clk_out
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__10074__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09220__A1 _04468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06034__A1 _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05468__S0 _01546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07782__A1 _03359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06585__A2 _02834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06952_ u_cpu.rf_ram.memory\[57\]\[5\] _03041_ _03047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09740_ _00194_ io_in[4] u_cpu.rf_ram.memory\[16\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
.ends

