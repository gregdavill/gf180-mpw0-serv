* NGSPICE file created from serv_2.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnq_1 D CLKN Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

.subckt serv_2 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_oeb[0] io_oeb[1] io_oeb[2]
+ io_oeb[3] io_oeb[4] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] vdd vss
XFILLER_95_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05903_ u_arbiter.i_wb_cpu_rdt\[22\] u_arbiter.i_wb_cpu_dbus_dat\[19\] _02431_ _02438_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09671_ _04638_ _04822_ _04830_ _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06883_ _02893_ _03079_ _03085_ _00378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06337__A2 _02756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07534__A1 _02717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05834_ _01444_ _02305_ _02393_ _02394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08622_ _04200_ _04211_ _00992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05640__S0 _01496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08553_ _03925_ _03974_ _04150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_05765_ _02336_ _02319_ _02338_ _02339_ _02340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_70_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07504_ u_cpu.rf_ram.memory\[134\]\[2\] _03435_ _03438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08484_ u_arbiter.i_wb_cpu_rdt\[24\] u_arbiter.i_wb_cpu_rdt\[8\] _02467_ _04088_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07837__A2 _03626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05696_ u_cpu.rf_ram.regzero _02273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_23_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07435_ _03314_ _03395_ _03399_ _00616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07366_ u_cpu.rf_ram.memory\[143\]\[5\] _03355_ _03361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09105_ u_cpu.rf_ram.memory\[101\]\[1\] _04503_ _04505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06317_ u_cpu.rf_ram.memory\[7\]\[4\] _02745_ _02750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08798__B1 _04311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05787__B _02292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08262__A2 _03885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07297_ _02666_ _03322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10417__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09036_ _04442_ _04463_ _04467_ _01150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06248_ _02669_ _02707_ _02708_ _00120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08014__A2 _03730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06179_ _02628_ _02657_ _02658_ _00101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05459__S0 _01529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10567__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06576__A2 _02900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07773__A1 _03508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09938_ _00332_ io_in[4] u_cpu.rf_ram.memory\[76\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09869_ _00263_ io_in[4] u_cpu.rf_ram.memory\[16\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07525__A1 _03314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06328__A2 _02756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05631__S0 _01551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09278__A1 _04448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07828__A2 _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10713_ _01083_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06500__A2 _02851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10644_ _01017_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10575_ _00948_ io_in[4] u_cpu.rf_ram.memory\[113\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10097__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09450__A1 _04638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08253__A2 _03885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09202__A1 _04444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08005__A2 _02954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11127_ _00058_ io_in[0] u_scanchain_local.module_data_in\[39\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11058_ _01426_ io_in[4] u_cpu.rf_ram.memory\[23\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06319__A2 _02745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07516__A1 _02675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10009_ _00403_ io_in[4] u_cpu.rf_ram.memory\[63\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05622__S0 _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05542__A3 _02101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05550_ _01566_ _02128_ _01480_ _02129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07819__A2 _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05481_ _01554_ _02060_ _01607_ _02061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08492__A2 _04024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07220_ _02803_ _02976_ _03276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07151_ _03098_ _03237_ _03238_ _00493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09732__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08244__A2 _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06102_ u_cpu.cpu.bufreg.c_r _02591_ _02592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_121_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07082_ u_cpu.rf_ram.memory\[56\]\[2\] _03197_ _03200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06033_ _02535_ _00078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__06007__A1 _02418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09882__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06558__A2 _02883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07755__A1 _03508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07984_ _03705_ _03710_ _03717_ _00848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09723_ _00117_ io_in[4] u_cpu.rf_ram.memory\[81\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06935_ _03098_ _03117_ _03118_ _00397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07507__A1 _03314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09654_ _02626_ _02838_ _04821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06866_ u_cpu.rf_ram.memory\[66\]\[6\] _03069_ _03076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08180__A1 u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08605_ _04186_ _04187_ _03912_ _04195_ _04196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_55_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05613__S0 _01495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05817_ _01467_ _02369_ _02382_ _00009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09585_ _04622_ _04782_ _04783_ _01383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06797_ _02618_ _02674_ _03037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06730__A2 _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08536_ u_cpu.cpu.immdec.imm30_25\[4\] _04102_ _04124_ u_cpu.cpu.immdec.imm30_25\[5\]
+ _04131_ _03959_ _04135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
X_05748_ u_cpu.cpu.state.o_cnt\[2\] _02291_ u_cpu.cpu.mem_bytecnt\[1\] _02323_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_23_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08467_ u_cpu.cpu.immdec.imm24_20\[2\] _04073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05679_ _02247_ _02256_ _02257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08483__A2 _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05297__A2 _01869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06494__A1 _02685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07418_ u_cpu.rf_ram.memory\[39\]\[4\] _03385_ _03390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08398_ _04011_ _04017_ _04018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07349_ _03318_ _03345_ _03351_ _00578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09432__A1 _04638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08235__A2 _03835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07288__I _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05310__B _01519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10360_ _00020_ io_in[4] u_cpu.rf_ram_if.rdata1\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06192__I _02631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07994__A1 _03697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09019_ u_cpu.rf_ram.memory\[95\]\[4\] _04453_ _04458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10291_ _00677_ io_in[4] u_cpu.rf_ram.memory\[130\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06920__I _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06549__A2 _02883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09499__A1 _04723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04980__A1 _01464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08171__A1 u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08171__B2 _02922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05604__S0 _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06721__A2 _02988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05080__S1 _01532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09755__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09671__A1 _04638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08474__A2 _03908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06485__A1 _02782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10732__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10627_ _01000_ io_in[4] u_cpu.rf_ram.memory\[32\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08226__A2 _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10558_ _00931_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06788__A2 _03028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10489_ _00862_ io_in[4] u_cpu.rf_ram.memory\[8\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05460__A2 _02039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10882__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07737__A1 _03508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08934__B1 _03909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10112__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04981_ _01504_ _01566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06960__A2 _03127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06720_ _02893_ _02988_ _02994_ _00306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08162__A1 u_arbiter.i_wb_cpu_dbus_dat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06651_ _02782_ _02954_ _02955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06712__A2 _02988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05602_ u_cpu.rf_ram.memory\[4\]\[7\] u_cpu.rf_ram.memory\[5\]\[7\] u_cpu.rf_ram.memory\[6\]\[7\]
+ u_cpu.rf_ram.memory\[7\]\[7\] _01523_ _01525_ _02180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10262__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05071__S1 _01509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09370_ _02647_ _04651_ _04655_ _01296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06582_ u_cpu.rf_ram.memory\[4\]\[7\] _02900_ _02908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_17_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08321_ _03906_ _03948_ _03949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05533_ _01543_ _02111_ _02112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08465__A2 _04069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08252_ u_cpu.rf_ram.memory\[113\]\[1\] _03885_ _03887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05464_ u_cpu.rf_ram.memory\[124\]\[5\] u_cpu.rf_ram.memory\[125\]\[5\] u_cpu.rf_ram.memory\[126\]\[5\]
+ u_cpu.rf_ram.memory\[127\]\[5\] _01496_ _01594_ _02044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_21_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07203_ _03266_ _03267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08183_ u_arbiter.i_wb_cpu_dbus_dat\[9\] _03835_ _03842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09414__A1 _04638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08217__A2 _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05395_ u_cpu.rf_ram.memory\[64\]\[4\] u_cpu.rf_ram.memory\[65\]\[4\] u_cpu.rf_ram.memory\[66\]\[4\]
+ u_cpu.rf_ram.memory\[67\]\[4\] _01522_ _01622_ _01976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_118_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07134_ u_cpu.rf_ram.memory\[53\]\[1\] _03227_ _03229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07976__A1 _03697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06779__A2 _02849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07065_ _03104_ _03187_ _03190_ _00455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06016_ u_cpu.cpu.ctrl.o_ibus_adr\[13\] u_cpu.cpu.ctrl.o_ibus_adr\[12\] _02499_ _02520_
+ _02521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_82_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05784__C _02265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08160__C _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05203__A2 _01785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07967_ u_cpu.rf_ram.memory\[120\]\[7\] _03693_ _03708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09706_ _00100_ io_in[4] u_cpu.rf_ram.memory\[82\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06918_ u_cpu.rf_ram.memory\[29\]\[3\] _03100_ _03107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10605__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04962__A1 _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07898_ _03502_ _03662_ _03666_ _00813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08153__A1 u_arbiter.i_wb_cpu_dbus_dat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09637_ _04811_ _04812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06849_ _02895_ _03059_ _03066_ _00363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09778__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06703__A2 _02978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07900__A1 _03504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05305__B _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09568_ u_cpu.rf_ram.memory\[25\]\[1\] _04772_ _04774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10755__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08519_ _03958_ _03929_ _04058_ _04119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_12_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05024__C _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09653__A1 _04638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08456__A2 _03941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09499_ _04723_ _04730_ _04731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_70_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08700__I0 u_arbiter.i_wb_cpu_dbus_adr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08208__A2 _03822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06219__A1 _02689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10412_ _00785_ io_in[4] u_cpu.rf_ram.memory\[91\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05690__A2 _02264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10343_ _00729_ io_in[4] u_cpu.rf_ram.memory\[125\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08351__B _03972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10274_ _00660_ io_in[4] u_cpu.rf_ram.memory\[133\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10135__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07719__A1 _03508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08392__A1 _03899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07195__A2 _03257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06942__A2 _03117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10285__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08144__A1 u_arbiter.i_wb_cpu_dbus_dat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06458__A1 _02687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05681__A2 u_cpu.cpu.state.o_cnt_r\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05180_ u_cpu.rf_ram.memory\[60\]\[2\] u_cpu.rf_ram.memory\[61\]\[2\] u_cpu.rf_ram.memory\[62\]\[2\]
+ u_cpu.rf_ram.memory\[63\]\[2\] _01562_ _01563_ _01763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_127_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05433__A2 _02012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06560__I _02661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11060__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08870_ u_cpu.rf_ram.memory\[109\]\[7\] _04351_ _04359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10628__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07186__A2 _03257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07821_ u_cpu.rf_ram.memory\[91\]\[2\] _03616_ _03619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09920__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05292__S1 _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04964_ u_cpu.rf_ram.memory\[32\]\[0\] u_cpu.rf_ram.memory\[33\]\[0\] u_cpu.rf_ram.memory\[34\]\[0\]
+ u_cpu.rf_ram.memory\[35\]\[0\] _01495_ _01499_ _01549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_42_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07752_ u_cpu.rf_ram.memory\[38\]\[5\] _03573_ _03579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08135__A1 u_arbiter.i_wb_cpu_dbus_dat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06703_ u_cpu.rf_ram.memory\[129\]\[6\] _02978_ _02985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10778__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07683_ _03508_ _03533_ _03540_ _00723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_04895_ _01481_ _01482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08686__A2 _04247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09422_ _04628_ _04681_ _04684_ _01319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05044__S1 _01500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05125__B _01600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06634_ u_cpu.rf_ram.memory\[17\]\[0\] _02945_ _02946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09353_ u_cpu.rf_ram.memory\[59\]\[4\] _04641_ _04646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08438__A2 _04041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09635__A1 _04638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06565_ _02897_ _02883_ _02898_ _00247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10008__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08304_ u_arbiter.i_wb_cpu_rdt\[8\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[8\]
+ _02466_ _03932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05516_ u_cpu.rf_ram.memory\[0\]\[6\] u_cpu.rf_ram.memory\[1\]\[6\] u_cpu.rf_ram.memory\[2\]\[6\]
+ u_cpu.rf_ram.memory\[3\]\[6\] _01508_ _01532_ _02095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09284_ _04434_ _04603_ _04604_ _01261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06496_ _02687_ _02851_ _02856_ _00220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07110__A2 _03207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05121__A1 _01490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08235_ _02445_ _03835_ _03876_ _00940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05447_ _01548_ _02026_ _01480_ _02027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05378_ u_cpu.rf_ram.memory\[120\]\[4\] u_cpu.rf_ram.memory\[121\]\[4\] u_cpu.rf_ram.memory\[122\]\[4\]
+ u_cpu.rf_ram.memory\[123\]\[4\] _01598_ _01556_ _01959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08166_ u_arbiter.i_wb_cpu_dbus_dat\[5\] _02915_ _03827_ _03829_ _03830_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__10158__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07117_ _03102_ _03217_ _03219_ _00478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08097_ u_cpu.rf_ram.memory\[116\]\[0\] _03780_ _03781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08610__A2 _04165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06621__A1 _02887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07048_ u_cpu.rf_ram.memory\[58\]\[3\] _03177_ _03181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07177__A2 _03247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08374__A1 _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08999_ _04444_ _04436_ _04445_ _01135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06924__A2 _03100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05283__S1 _01500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04935__A1 _01506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08126__A1 _03703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10961_ _01330_ io_in[4] u_cpu.rf_ram.memory\[111\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06137__B1 u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08677__A2 _04247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06688__A1 _02608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10892_ _01261_ io_in[4] u_cpu.rf_ram.memory\[108\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08429__A2 _04041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04874__B u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07101__A2 _03207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11083__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06612__A1 _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05415__A2 _01995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10326_ _00712_ io_in[4] u_cpu.rf_ram.memory\[127\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_4_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09943__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10257_ _00643_ io_in[4] u_cpu.rf_ram.memory\[135\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07168__A2 _03247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08365__A1 _03974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10188_ _00574_ io_in[4] u_cpu.rf_ram.memory\[70\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05179__B2 _01761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06915__A2 _03100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05718__A3 _02292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10920__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05274__S1 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04926__A1 _01506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08668__A2 _04237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06679__A1 _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05026__S1 _01563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07340__A2 _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09617__A1 _02693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06350_ u_cpu.rf_ram.memory\[78\]\[0\] _02770_ _02771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05301_ _01597_ _01882_ _01600_ _01883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10300__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06281_ u_cpu.rf_ram.memory\[20\]\[7\] _02719_ _02727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08840__A2 _04327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05232_ u_cpu.rf_ram.memory\[140\]\[2\] u_cpu.rf_ram.memory\[141\]\[2\] u_cpu.rf_ram.memory\[142\]\[2\]
+ u_cpu.rf_ram.memory\[143\]\[2\] _01634_ _01635_ _01815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08020_ _02662_ _03730_ _03737_ _00864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06851__A1 _02897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05163_ _01493_ _01745_ _01746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10450__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06603__A1 _02305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09971_ _00365_ io_in[4] u_cpu.rf_ram.memory\[66\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05094_ u_cpu.rf_ram.memory\[56\]\[1\] u_cpu.rf_ram.memory\[57\]\[1\] u_cpu.rf_ram.memory\[58\]\[1\]
+ u_cpu.rf_ram.memory\[59\]\[1\] _01567_ _01568_ _01678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_115_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08922_ u_cpu.rf_ram.memory\[93\]\[6\] _04381_ _04388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08356__A1 _03914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07159__A2 _03237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08853_ u_cpu.cpu.immdec.imm11_7\[2\] _02624_ _02729_ _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_112_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07804_ _02395_ _03608_ _00776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05265__S1 _01531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08784_ u_arbiter.i_wb_cpu_ibus_adr\[0\] _04309_ _04311_ u_arbiter.i_wb_cpu_ibus_adr\[1\]
+ _04312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_73_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08108__A1 _03703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05996_ _02389_ u_scanchain_local.module_data_in\[49\] _02506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07735_ _03506_ _03563_ _03569_ _00746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04947_ _01531_ _01532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08659__A2 _04237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07666_ u_cpu.rf_ram.memory\[127\]\[7\] _03523_ _03531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04878_ _01464_ _01465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_129_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07331__A2 _03335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09405_ u_cpu.rf_ram.memory\[110\]\[3\] _04671_ _04675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06617_ _02881_ _02935_ _02936_ _00261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09608__A1 u_cpu.rf_ram.memory\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07597_ _02647_ _03485_ _03489_ _00688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09336_ _04634_ _04624_ _04635_ _01282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09816__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06548_ _02641_ _02887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09267_ u_cpu.rf_ram.memory\[83\]\[1\] _04593_ _04595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06479_ _02689_ _02840_ _02846_ _00213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05645__A2 _02222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08218_ _03864_ _03865_ _00934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09198_ _04440_ _04553_ _04556_ _01223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09966__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08149_ _03815_ _00915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_88_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08595__A1 _03909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07398__A2 _03375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11160_ io_oeb[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_106_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10943__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10111_ _00505_ io_in[4] u_cpu.rf_ram.memory\[9\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11091_ _00059_ io_in[0] u_arbiter.i_wb_cpu_rdt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10042_ _00436_ io_in[4] u_cpu.rf_ram.memory\[19\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08898__A2 _04371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05256__S1 _01532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07570__A2 _02976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05581__A1 _02140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10944_ _01313_ io_in[4] u_cpu.rf_ram.memory\[110\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06125__A3 _02606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07322__A2 _03335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10323__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10875_ _01244_ io_in[4] u_cpu.rf_ram.memory\[106\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08822__A2 _04327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10473__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05636__A2 _02213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06833__A1 _02897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08586__A1 _03986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07389__A2 _03365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10309_ _00695_ io_in[4] u_cpu.rf_ram.memory\[22\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08338__A1 _03904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08889__A2 _04361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05247__S1 _01509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07010__A1 u_cpu.rf_ram.memory\[19\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05850_ u_cpu.cpu.bne_or_bge _02306_ _02407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07561__A2 _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05572__A1 _01621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05781_ u_arbiter.i_wb_cpu_dbus_dat\[0\] u_arbiter.i_wb_cpu_dbus_dat\[8\] u_arbiter.i_wb_cpu_dbus_dat\[16\]
+ u_arbiter.i_wb_cpu_dbus_dat\[24\] _02306_ _02355_ _02356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_81_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07520_ u_cpu.rf_ram.memory\[133\]\[1\] _03445_ _03447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09839__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08510__A1 _03932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07313__A2 _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07451_ _03312_ _03405_ _03408_ _00623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_63_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06402_ u_cpu.rf_ram.memory\[46\]\[6\] _02794_ _02801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10816__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07382_ u_cpu.rf_ram.memory\[14\]\[4\] _03365_ _03370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09066__A2 _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09121_ u_cpu.rf_ram.memory\[102\]\[0\] _04513_ _04514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06333_ _02683_ _02756_ _02759_ _00154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09989__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09052_ u_cpu.rf_ram.memory\[28\]\[0\] _04476_ _04477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06264_ _02674_ _02716_ _02717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05478__I2 u_cpu.rf_ram.memory\[82\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08003_ u_cpu.rf_ram.memory\[121\]\[7\] _03720_ _03728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05215_ _01602_ _01797_ _01798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10966__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06195_ _02617_ _02671_ _02672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__08577__B2 _04003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05146_ u_cpu.rf_ram.memory\[136\]\[1\] u_cpu.rf_ram.memory\[137\]\[1\] u_cpu.rf_ram.memory\[138\]\[1\]
+ u_cpu.rf_ram.memory\[139\]\[1\] _01641_ _01642_ _01730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_104_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09954_ _00348_ io_in[4] u_cpu.rf_ram.memory\[6\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05077_ _01528_ _01660_ _01534_ _01661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_44_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08905_ _02662_ _04371_ _04378_ _01108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09885_ _00279_ io_in[4] u_cpu.rf_ram.memory\[40\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07001__A1 _03112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08836_ u_cpu.cpu.ctrl.o_ibus_adr\[25\] _04327_ _04329_ u_cpu.cpu.ctrl.o_ibus_adr\[26\]
+ _04339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07552__A2 _02976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10346__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05563__A1 _01464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08767_ _03695_ _04299_ _04301_ _01047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05979_ u_cpu.cpu.ctrl.o_ibus_adr\[9\] _02492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_26_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07718_ u_cpu.rf_ram.memory\[124\]\[6\] _03553_ _03560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08698_ u_arbiter.i_wb_cpu_dbus_adr\[6\] u_arbiter.i_wb_cpu_dbus_adr\[7\] _04257_
+ _04262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_25_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08501__A1 _03955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07304__A2 _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07649_ _03510_ _03513_ _03521_ _00708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10496__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10660_ _01033_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05410__S1 _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09057__A2 _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09319_ _04623_ _04624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_139_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08804__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10591_ _00964_ io_in[4] u_cpu.cpu.decode.op22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08624__B _04013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06815__A1 _02667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06923__I _02656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06291__A2 _02733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08568__A1 _02259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11143_ _00076_ io_in[0] u_scanchain_local.module_data_in\[55\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11121__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07791__A2 _03593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11074_ _01434_ io_in[4] u_cpu.rf_ram_if.rgnt vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10025_ _00419_ io_in[4] u_cpu.rf_ram.memory\[61\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07543__A2 _03455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10839__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09296__A2 _04603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10927_ _01296_ io_in[4] u_cpu.rf_ram.memory\[10\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05401__S1 _01500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05857__A2 _02355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10858_ _01227_ io_in[4] u_cpu.rf_ram.memory\[79\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10989__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10789_ _01158_ io_in[4] u_cpu.rf_ram.memory\[28\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05609__A2 _02186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06282__A2 _02719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10219__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05000_ u_cpu.rf_ram.memory\[100\]\[0\] u_cpu.rf_ram.memory\[101\]\[0\] u_cpu.rf_ram.memory\[102\]\[0\]
+ u_cpu.rf_ram.memory\[103\]\[0\] _01572_ _01573_ _01585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_67_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08559__B2 _03914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09220__A2 _04563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07231__A1 _03108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05468__S1 _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07782__A2 _03593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10369__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06951_ _03126_ _03127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05793__A1 _02305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05902_ _02437_ _00042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_41_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09670_ u_cpu.rf_ram.memory\[89\]\[7\] _04822_ _04830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06882_ u_cpu.rf_ram.memory\[65\]\[5\] _03079_ _03085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08696__S _04257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07534__A2 _02976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08621_ _03959_ _04202_ _04208_ _04210_ _04211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_39_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05833_ u_cpu.cpu.state.init_done _02392_ _02393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__04979__S0 _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08552_ _03969_ _04148_ _04149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05640__S1 _01594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05764_ u_cpu.cpu.ctrl.pc_plus_offset_cy_r _02330_ _02339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09287__A2 _04603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07503_ _03310_ _03435_ _03437_ _00646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08483_ _03922_ _03918_ _04086_ _03940_ _04023_ _04087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_35_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05695_ u_cpu.rf_ram_if.rtrig1 _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05848__A2 _02389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07434_ u_cpu.rf_ram.memory\[137\]\[3\] _03395_ _03399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09039__A2 _04463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07365_ _03316_ _03355_ _03360_ _00585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08444__B _03915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09104_ _04434_ _04503_ _04504_ _01181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08798__A1 u_cpu.cpu.ctrl.o_ibus_adr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06316_ _02647_ _02745_ _02749_ _00147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07296_ _03320_ _03308_ _03321_ _00555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09035_ u_cpu.rf_ram.memory\[96\]\[3\] _04463_ _04467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06273__A2 _02719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06247_ u_cpu.rf_ram.memory\[18\]\[0\] _02707_ _02708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11144__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06178_ u_cpu.rf_ram.memory\[82\]\[5\] _02628_ _02658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09211__A2 _04563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05459__S1 _01500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05129_ _01617_ _01712_ _01607_ _01713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_85_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08970__A1 _03695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07773__A2 _03583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09937_ _00331_ io_in[4] u_cpu.rf_ram.memory\[76\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05784__A1 _01442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09868_ _00262_ io_in[4] u_cpu.rf_ram.memory\[16\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07525__A2 _03445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08819_ _04330_ _01070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09799_ _00193_ io_in[4] u_cpu.rf_ram.memory\[44\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05631__S1 _01524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09278__A2 _04593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10712_ _01082_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05395__S0 _01522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10643_ _01016_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10574_ _00947_ io_in[4] u_cpu.rf_ram.memory\[113\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09450__A2 _04691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07461__A1 _03322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09202__A2 _04553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10511__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07213__A1 _03108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08961__A1 _03965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07764__A2 _03583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11126_ _00057_ io_in[0] u_scanchain_local.module_data_in\[38\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05775__A1 _01443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05775__B2 _02334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11057_ _01425_ io_in[4] u_cpu.rf_ram.memory\[23\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10661__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07516__A2 _02976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10008_ _00402_ io_in[4] u_cpu.rf_ram.memory\[63\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08529__B _04052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05622__S1 _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09269__A2 _04593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11017__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05480_ u_cpu.rf_ram.memory\[84\]\[5\] u_cpu.rf_ram.memory\[85\]\[5\] u_cpu.rf_ram.memory\[86\]\[5\]
+ u_cpu.rf_ram.memory\[87\]\[5\] _01507_ _01605_ _02060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__05386__S0 _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08229__B1 _03808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10041__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07150_ u_cpu.rf_ram.memory\[52\]\[0\] _03237_ _03238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06563__I _02666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09441__A2 _04691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06101_ u_cpu.cpu.alu.i_rs1 _02584_ _02585_ _02591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_34_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06255__A2 _02707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07452__A1 u_cpu.rf_ram.memory\[49\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07081_ _03102_ _03197_ _03199_ _00462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06032_ _02389_ u_scanchain_local.module_data_in\[56\] _02534_ _02535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10191__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08952__A1 u_cpu.cpu.immdec.imm11_7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07755__A2 _03573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07983_ u_cpu.rf_ram.memory\[118\]\[6\] _03710_ _03717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09722_ _00116_ io_in[4] u_cpu.rf_ram.memory\[81\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06934_ u_cpu.rf_ram.memory\[63\]\[0\] _03117_ _03118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07507__A2 _03435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09653_ _04638_ _04812_ _04820_ _01414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06865_ _02893_ _03069_ _03075_ _00370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08604_ _04192_ _04193_ _04194_ _04195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__08180__A2 _03835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05816_ u_cpu.rf_ram_if.rdata0\[2\] _01467_ _02382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09584_ u_cpu.rf_ram.memory\[24\]\[0\] _04782_ _04783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05613__S1 _01499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06191__A1 _02628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06796_ _02897_ _03028_ _03036_ _00340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_70_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08535_ _03966_ _04130_ _04133_ _04134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_82_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05747_ _02263_ _02320_ _02321_ _02322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_70_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08466_ _04029_ _04072_ _00975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05678_ _02249_ _02251_ _02253_ _02255_ _01466_ _02256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__09680__A2 _04832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07417_ _03314_ _03385_ _03389_ _00608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05297__A3 _01878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06494__A2 _02851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07691__A1 _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08397_ _02911_ _03904_ _04014_ _04016_ _04017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_137_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07348_ u_cpu.rf_ram.memory\[70\]\[5\] _03345_ _03351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09432__A2 _04681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10534__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07443__A1 _03322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07279_ _02636_ _03310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07994__A2 _03720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09018_ _04442_ _04453_ _04457_ _01142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10290_ _00676_ io_in[4] u_cpu.rf_ram.memory\[131\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09196__A1 _04438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10684__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08943__A1 _03924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07746__A2 _03573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04980__A2 _01564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08171__A2 _03808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05604__S1 _01509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10064__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09671__A2 _04822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06485__A2 _02849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05501__B _01482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10626_ _00999_ io_in[4] u_cpu.rf_ram.memory\[32\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09423__A2 _04681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06237__A2 _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10557_ _00930_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07985__A2 _03710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08304__S _02466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10488_ _00861_ io_in[4] u_cpu.rf_ram.memory\[8\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05996__A1 _02389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07737__A2 _03563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08934__A1 _03944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08934__B2 _03932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11109_ _00039_ io_in[0] u_arbiter.i_wb_cpu_rdt\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_04980_ _01464_ _01564_ _01565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10407__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06650_ _02716_ _02779_ _02954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_65_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06173__A1 _02628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05601_ _02172_ _02174_ _02176_ _02178_ _01486_ _02179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_92_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06581_ _02662_ _02900_ _02907_ _00254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_45_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08320_ _03946_ _03947_ _03948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05532_ u_cpu.rf_ram.memory\[60\]\[6\] u_cpu.rf_ram.memory\[61\]\[6\] u_cpu.rf_ram.memory\[62\]\[6\]
+ u_cpu.rf_ram.memory\[63\]\[6\] _01496_ _01594_ _02111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_33_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09662__A2 _04822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10557__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08251_ _03691_ _03885_ _03886_ _00946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06476__A2 _02840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05463_ _02036_ _02038_ _02040_ _02042_ _01560_ _02043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__07673__A1 _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07202_ _02766_ _02976_ _03266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08182_ _03840_ _03841_ _00922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05394_ _01968_ _01970_ _01972_ _01974_ _01486_ _01975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__09414__A2 _04671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07133_ _03098_ _03227_ _03228_ _00485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07425__A1 _03322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05130__C _01486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07976__A2 _03710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07064_ u_cpu.rf_ram.memory\[57\]\[2\] _03187_ _03190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09178__A1 _04438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06015_ u_cpu.cpu.ctrl.o_ibus_adr\[17\] u_cpu.cpu.ctrl.o_ibus_adr\[16\] u_cpu.cpu.ctrl.o_ibus_adr\[15\]
+ u_cpu.cpu.ctrl.o_ibus_adr\[14\] _02520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_47_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07728__A2 _03563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08925__A1 _03707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05739__A1 _02313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06400__A2 _02794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07966_ _02666_ _03707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09705_ _00099_ io_in[4] u_cpu.rf_ram.memory\[82\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_101_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06917_ _02646_ _03106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07897_ u_cpu.rf_ram.memory\[35\]\[3\] _03662_ _03666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10087__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09350__A1 _04628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09636_ _02717_ _04349_ _04811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06848_ u_cpu.rf_ram.memory\[67\]\[6\] _03059_ _03066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07900__A2 _03662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09567_ _04622_ _04772_ _04773_ _01375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06779_ _02768_ _02849_ _03027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08518_ _03924_ _03918_ _03988_ _04000_ _04118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_54_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09498_ _02305_ _02400_ _04729_ u_cpu.cpu.state.genblk1.misalign_trap_sync_r _04726_
+ _04730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__09653__A2 _04812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08449_ _04000_ _03929_ _03975_ _03972_ _04058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_11_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05321__B _01482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09405__A2 _04671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06219__A2 _02679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10411_ _00784_ io_in[4] u_cpu.rf_ram.memory\[91\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07967__A2 _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10342_ _00728_ io_in[4] u_cpu.rf_ram.memory\[125\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08351__C _03975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10273_ _00659_ io_in[4] u_cpu.rf_ram.memory\[133\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07719__A2 _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08392__A2 _03917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09722__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08144__A2 u_arbiter.i_wb_cpu_dbus_dat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06155__A1 _02628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09872__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09644__A2 _04812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07655__A1 _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06458__A2 _02829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05130__A2 _01709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10609_ _00982_ io_in[4] u_cpu.cpu.immdec.imm30_25\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07407__A1 _03322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05681__A3 u_cpu.cpu.state.o_cnt_r\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07958__A2 _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08080__A1 _03691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05969__A1 u_cpu.cpu.ctrl.o_ibus_adr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06630__A2 _02935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08907__A1 _02667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07820_ _03498_ _03616_ _03618_ _00782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07751_ _03504_ _03573_ _03578_ _00753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_04963_ _01504_ _01548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_77_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08135__A2 _02915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06702_ _02893_ _02978_ _02984_ _00298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_93_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07682_ u_cpu.rf_ram.memory\[126\]\[6\] _03533_ _03540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04894_ _01480_ _01481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09421_ u_cpu.rf_ram.memory\[86\]\[2\] _04681_ _04684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06633_ _02944_ _02945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06697__A2 _02978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07894__A1 _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09352_ _04630_ _04641_ _04645_ _01288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06564_ u_cpu.rf_ram.memory\[50\]\[7\] _02883_ _02898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09635__A2 _04802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08303_ _03918_ _03930_ _03931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_100_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05515_ _01493_ _02093_ _02094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06449__A2 _02829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07646__A1 u_cpu.rf_ram.memory\[128\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09283_ u_cpu.rf_ram.memory\[108\]\[0\] _04603_ _04604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06495_ u_cpu.rf_ram.memory\[43\]\[4\] _02851_ _02856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05141__B _01471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08234_ u_arbiter.i_wb_cpu_rdt\[26\] _02924_ _03874_ u_arbiter.i_wb_cpu_dbus_dat\[27\]
+ _03876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_21_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05446_ u_cpu.rf_ram.memory\[56\]\[5\] u_cpu.rf_ram.memory\[57\]\[5\] u_cpu.rf_ram.memory\[58\]\[5\]
+ u_cpu.rf_ram.memory\[59\]\[5\] _01567_ _01568_ _02026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__05121__A2 _01695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08165_ _03828_ _03829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05377_ _01543_ _01957_ _01958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07949__A2 _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07116_ u_cpu.rf_ram.memory\[54\]\[1\] _03217_ _03219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08096_ _03779_ _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_106_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06082__B1 _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06621__A2 _02935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07047_ _03104_ _03177_ _03180_ _00447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09745__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09571__A1 _04628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08374__A2 u_arbiter.i_wb_cpu_rdt\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08998_ u_cpu.rf_ram.memory\[94\]\[4\] _04436_ _04445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05188__A2 _01766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06385__A1 _02691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07949_ u_cpu.rf_ram.memory\[120\]\[1\] _03693_ _03696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04935__A2 _01516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10722__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08126__A2 _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10960_ _01329_ io_in[4] u_cpu.rf_ram.memory\[111\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06137__A1 _02606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09895__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09503__S _04723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09619_ _04801_ _04802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06688__A2 _02622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05035__C _01486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10891_ _01260_ io_in[4] u_cpu.rf_ram.memory\[83\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06926__I _02661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10872__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09626__A2 _04802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04874__C _01460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07637__A1 _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08834__B1 _04329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10102__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06860__A2 _03069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08062__A1 _03691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10325_ _00711_ io_in[4] u_cpu.rf_ram.memory\[127\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10252__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10256_ _00642_ io_in[4] u_cpu.rf_ram.memory\[135\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08365__A2 _03908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10187_ _00573_ io_in[4] u_cpu.rf_ram.memory\[70\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05179__A2 _01757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05718__A4 _02293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04926__A2 _01510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09314__A1 _04448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08117__A2 _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05226__B _01481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06128__A1 _01460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07876__A1 _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06679__A2 _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09617__A2 _04792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07628__A1 _03508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05300_ u_cpu.rf_ram.memory\[88\]\[3\] u_cpu.rf_ram.memory\[89\]\[3\] u_cpu.rf_ram.memory\[90\]\[3\]
+ u_cpu.rf_ram.memory\[91\]\[3\] _01598_ _01556_ _01882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_72_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06280_ _02691_ _02719_ _02726_ _00134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06300__A1 _02657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05231_ _01465_ _01813_ _01814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06851__A2 _03059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05162_ u_cpu.rf_ram.memory\[4\]\[2\] u_cpu.rf_ram.memory\[5\]\[2\] u_cpu.rf_ram.memory\[6\]\[2\]
+ u_cpu.rf_ram.memory\[7\]\[2\] _01523_ _01525_ _01745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_144_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09768__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09970_ _00364_ io_in[4] u_cpu.rf_ram.memory\[67\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07800__A1 _02291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05093_ _01464_ _01676_ _01677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08921_ _03703_ _04381_ _04387_ _01115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10745__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09553__A1 _04628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08356__A2 _03908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08852_ _04348_ _01085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_111_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07803_ u_cpu.cpu.mem_bytecnt\[1\] _03607_ _03608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08783_ _04310_ _04311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05995_ u_arbiter.i_wb_cpu_dbus_adr\[12\] _02397_ _02504_ _02505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08108__A2 _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07734_ u_cpu.rf_ram.memory\[123\]\[5\] _03563_ _03569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04946_ _01498_ _01531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06119__A1 u_cpu.cpu.immdec.imm11_7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10895__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07665_ _03508_ _03523_ _03530_ _00715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07867__A1 u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04877_ _01463_ _01464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09404_ _04628_ _04671_ _04674_ _01311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06616_ u_cpu.rf_ram.memory\[16\]\[0\] _02935_ _02936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07596_ u_cpu.rf_ram.memory\[12\]\[3\] _03485_ _03489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_41_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09608__A2 _04792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10125__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09335_ u_cpu.rf_ram.memory\[84\]\[5\] _04624_ _04635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07619__A1 _03502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08166__C _03829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06547_ _02885_ _02883_ _02886_ _00241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09266_ _04434_ _04593_ _04594_ _01253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06478_ u_cpu.rf_ram.memory\[41\]\[5\] _02840_ _02846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08217_ u_arbiter.i_wb_cpu_rdt\[20\] _03807_ _03829_ u_arbiter.i_wb_cpu_dbus_dat\[21\]
+ _03865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05429_ _01528_ _02008_ _01534_ _02009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09197_ u_cpu.rf_ram.memory\[79\]\[2\] _04553_ _04556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06842__A2 _03059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10275__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08044__A1 _03691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08148_ u_arbiter.i_wb_cpu_rdt\[1\] _02924_ _03814_ _03815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08079_ u_cpu.rf_ram.memory\[115\]\[0\] _03770_ _03771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10110_ _00504_ io_in[4] u_cpu.rf_ram.memory\[9\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11090_ _00048_ io_in[0] u_arbiter.i_wb_cpu_rdt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10041_ _00435_ io_in[4] u_cpu.rf_ram.memory\[19\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10943_ _01312_ io_in[4] u_cpu.rf_ram.memory\[110\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10874_ _01243_ io_in[4] u_cpu.rf_ram.memory\[106\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11050__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10618__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07086__A2 _03197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08283__A1 _03909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05097__A1 _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06833__A2 _03049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09910__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09083__I0 u_arbiter.i_wb_cpu_rdt\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10768__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08586__A2 _03906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06597__A1 u_arbiter.i_wb_cpu_dbus_dat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10308_ _00694_ io_in[4] u_cpu.rf_ram.memory\[22\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08312__S _02465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09535__A1 _04628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10239_ _00625_ io_in[4] u_cpu.rf_ram.memory\[49\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07010__A2 _03157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05780_ u_cpu.cpu.bufreg.lsb\[1\] _02355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05572__A2 _02150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10148__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08510__A2 _03988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07450_ u_cpu.rf_ram.memory\[49\]\[2\] _03405_ _03408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06401_ _02689_ _02794_ _02800_ _00181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07381_ _02647_ _03365_ _03369_ _00592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_34_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05403__C _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10298__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09120_ _04512_ _04513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06332_ u_cpu.rf_ram.memory\[80\]\[2\] _02756_ _02759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08274__A1 _02465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05088__A1 _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09051_ _04475_ _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06824__A2 _03049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06263_ _01563_ _02616_ _02716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_124_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08002_ _03705_ _03720_ _03727_ _00856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05214_ u_cpu.rf_ram.memory\[80\]\[2\] u_cpu.rf_ram.memory\[81\]\[2\] u_cpu.rf_ram.memory\[82\]\[2\]
+ u_cpu.rf_ram.memory\[83\]\[2\] _01544_ _01594_ _01797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_116_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08026__A1 _02632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06194_ _01498_ _02670_ _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_144_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08577__A2 _04165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05145_ _01638_ _01728_ _01482_ _01729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06588__A1 _02395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09953_ _00347_ io_in[4] u_cpu.rf_ram.memory\[6\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05076_ u_cpu.rf_ram.memory\[0\]\[1\] u_cpu.rf_ram.memory\[1\]\[1\] u_cpu.rf_ram.memory\[2\]\[1\]
+ u_cpu.rf_ram.memory\[3\]\[1\] _01530_ _01532_ _01660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_103_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05260__A1 _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09526__A1 u_cpu.cpu.genblk3.csr.o_new_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08904_ u_cpu.rf_ram.memory\[2\]\[6\] _04371_ _04378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09884_ _00278_ io_in[4] u_cpu.rf_ram.memory\[40\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07001__A2 _03147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08835_ _04338_ _01078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08766_ u_cpu.rf_ram.memory\[30\]\[1\] _04299_ _04301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05978_ _02488_ _02490_ _02491_ _00066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05563__A2 _02141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06760__A1 _02897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07717_ _03506_ _03553_ _03559_ _00738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11073__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04929_ u_cpu.rf_ram.memory\[20\]\[0\] u_cpu.rf_ram.memory\[21\]\[0\] u_cpu.rf_ram.memory\[22\]\[0\]
+ u_cpu.rf_ram.memory\[23\]\[0\] _01497_ _01501_ _01514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_2739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08697_ _04261_ _01017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08501__A2 _04101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07648_ u_cpu.rf_ram.memory\[128\]\[7\] _03513_ _03521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06512__A1 _02685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07579_ _03314_ _03475_ _03479_ _00680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09933__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09318_ _02626_ _02717_ _04623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08265__A1 _03707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07068__A2 _03187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10590_ _00963_ io_in[4] u_cpu.cpu.decode.op21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05079__A1 _01528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09249_ u_cpu.rf_ram.memory\[107\]\[1\] _04583_ _04585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10910__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06815__A2 _03039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05874__I0 u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06579__A1 _02657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11142_ _00075_ io_in[0] u_scanchain_local.module_data_in\[54\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07240__A2 _03287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05251__A1 _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09517__A1 _02301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11073_ _01433_ io_in[4] u_cpu.rf_ram_if.rdata0\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10024_ _00418_ io_in[4] u_cpu.rf_ram.memory\[61\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05003__A1 _01548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10440__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10926_ _01295_ io_in[4] u_cpu.rf_ram.memory\[10\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05306__A2 _01883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06503__A1 _02754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10857_ _01226_ io_in[4] u_cpu.rf_ram.memory\[79\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10788_ _01157_ io_in[4] u_cpu.rf_ram.memory\[28\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10590__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06806__A2 _03039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08008__A1 _02632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05490__A1 _01617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07231__A2 _03277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05242__A1 _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09508__A1 _02263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06950_ _02766_ _02827_ _03126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05793__A2 _02318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05901_ u_arbiter.i_wb_cpu_rdt\[21\] u_arbiter.i_wb_cpu_dbus_dat\[18\] _02431_ _02437_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09806__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11096__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06881_ _02891_ _03079_ _03084_ _00377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08620_ _04164_ _04209_ _04210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05832_ u_cpu.cpu.state.o_cnt_r\[1\] u_cpu.cpu.state.o_cnt_r\[0\] u_cpu.cpu.state.o_cnt_r\[3\]
+ u_cpu.cpu.state.o_cnt_r\[2\] _02392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_67_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06742__A1 _02897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04979__S1 _01563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08551_ _03925_ _04052_ _04148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05763_ _02319_ _02337_ _02338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09956__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07502_ u_cpu.rf_ram.memory\[134\]\[1\] _03435_ _03437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08482_ _03978_ _04086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_36_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07298__A2 _03308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05694_ _02263_ _02267_ _02268_ _02270_ _02271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_50_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07433_ _03312_ _03395_ _03398_ _00615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10933__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07364_ u_cpu.rf_ram.memory\[143\]\[4\] _03355_ _03360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09103_ u_cpu.rf_ram.memory\[101\]\[0\] _04503_ _04504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06315_ u_cpu.rf_ram.memory\[7\]\[3\] _02745_ _02749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08798__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07295_ u_cpu.rf_ram.memory\[72\]\[6\] _03308_ _03321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09034_ _04440_ _04463_ _04466_ _01149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06246_ _02706_ _02707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07470__A2 _03415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05481__A1 _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06177_ _02656_ _02657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08460__B _02259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05128_ u_cpu.rf_ram.memory\[84\]\[1\] u_cpu.rf_ram.memory\[85\]\[1\] u_cpu.rf_ram.memory\[86\]\[1\]
+ u_cpu.rf_ram.memory\[87\]\[1\] _01507_ _01605_ _01712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_116_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07222__A2 _03277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10313__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05233__A1 _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08970__A2 _04425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09936_ _00330_ io_in[4] u_cpu.rf_ram.memory\[76\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05059_ _01465_ _01643_ _01644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_131_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06981__A1 _03110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09867_ _00261_ io_in[4] u_cpu.rf_ram.memory\[16\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10463__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08818_ u_cpu.cpu.ctrl.o_ibus_adr\[16\] _04327_ _04329_ u_cpu.cpu.ctrl.o_ibus_adr\[17\]
+ _04330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_86_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09798_ _00192_ io_in[4] u_cpu.rf_ram.memory\[44\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05092__S0 _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08749_ _02590_ _02592_ _04287_ _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08486__A1 _03914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07289__A2 _03308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10711_ _01081_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05395__S1 _01622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10642_ _01015_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10573_ _00946_ io_in[4] u_cpu.rf_ram.memory\[113\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07461__A2 _03405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09829__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06016__A3 _02499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08410__A1 _04009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07213__A2 _03267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08410__B2 _03955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05224__A1 _01621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11125_ _00056_ io_in[0] u_scanchain_local.module_data_in\[37\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08961__A2 _03962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10806__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11056_ _01424_ io_in[4] u_cpu.rf_ram.memory\[23\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05218__C _01486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09979__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10007_ _00401_ io_in[4] u_cpu.rf_ram.memory\[63\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06724__A1 _02897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05083__S0 _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10956__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08477__A1 _04031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10909_ _01278_ io_in[4] u_cpu.rf_ram.memory\[84\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05386__S1 _01563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08229__A1 u_arbiter.i_wb_cpu_rdt\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08229__B2 u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06100_ _02322_ _02589_ _02590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07080_ u_cpu.rf_ram.memory\[56\]\[1\] _03197_ _03199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07452__A2 _03405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10336__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06031_ _02388_ _02532_ _02533_ _02534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_114_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07204__A2 _03267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05215__A1 _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08952__A2 _02392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07982_ _03703_ _03710_ _03716_ _00847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10486__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05409__B _01534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05766__A2 _02334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06963__A1 _03110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06933_ _03116_ _03117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09721_ _00115_ io_in[4] u_cpu.rf_ram.memory\[81\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09652_ u_cpu.rf_ram.memory\[100\]\[7\] _04812_ _04820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06864_ u_cpu.rf_ram.memory\[66\]\[5\] _03069_ _03075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06715__A1 u_cpu.rf_ram.memory\[139\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05074__S0 _01523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08603_ _04031_ _03961_ _04194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05815_ _01467_ _02274_ _02381_ _00008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09583_ _04781_ _04782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_43_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06795_ u_cpu.rf_ram.memory\[75\]\[7\] _03028_ _03036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06191__A2 _02667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08534_ _03906_ _04132_ _04133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08468__A1 u_cpu.cpu.immdec.imm24_20\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05746_ _02263_ _02267_ _02268_ _02321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_24_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08465_ u_cpu.cpu.immdec.imm24_20\[1\] _04069_ _04070_ u_cpu.cpu.immdec.imm24_20\[2\]
+ _04072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_23_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05677_ _01465_ _02254_ _01534_ _02255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07416_ u_cpu.rf_ram.memory\[39\]\[3\] _03385_ _03389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11111__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08396_ _03910_ _04015_ _04016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07691__A2 _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07347_ _03316_ _03345_ _03350_ _00577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08640__A1 _02305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07443__A2 _03395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07278_ _03306_ _03308_ _03309_ _00549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09017_ u_cpu.rf_ram.memory\[95\]\[3\] _04453_ _04457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05454__A1 _01492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06229_ u_cpu.rf_ram.memory\[81\]\[0\] _02697_ _02698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10829__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09196__A2 _04553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09919_ _00313_ io_in[4] u_cpu.rf_ram.memory\[77\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10979__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06929__I _02666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06706__A1 _02897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05065__S0 _01497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10209__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07682__A2 _03533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10359__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05693__A1 _02263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10625_ _00998_ io_in[4] u_cpu.rf_ram.memory\[32\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10556_ _00929_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07434__A2 _03395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05445__A1 _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10487_ _00860_ io_in[4] u_cpu.rf_ram.memory\[8\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09187__A2 _04543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04912__I _01496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05229__B _01471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08934__A2 _03908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05748__A2 _02291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06945__A1 _03110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11108_ _00038_ io_in[0] u_arbiter.i_wb_cpu_rdt\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11039_ _01408_ io_in[4] u_cpu.rf_ram.memory\[100\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06173__A2 _02652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05600_ _01506_ _02177_ _01519_ _02178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_24_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11134__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06580_ u_cpu.rf_ram.memory\[4\]\[6\] _02900_ _02907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09111__A2 _04503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05531_ _02103_ _02105_ _02107_ _02109_ _01560_ _02110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_127_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08250_ u_cpu.rf_ram.memory\[113\]\[0\] _03885_ _03886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05462_ _01566_ _02041_ _01558_ _02042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07673__A2 _03533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07201_ _02667_ _03257_ _03265_ _00516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05684__A1 u_arbiter.i_wb_cpu_dbus_we vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08181_ u_arbiter.i_wb_cpu_rdt\[8\] _03822_ _03833_ u_arbiter.i_wb_cpu_dbus_dat\[9\]
+ _03841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05393_ _01554_ _01973_ _01607_ _01974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07132_ u_cpu.rf_ram.memory\[53\]\[0\] _03227_ _03228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07425__A2 _03385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05436__A1 _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07063_ _03102_ _03187_ _03189_ _00454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06014_ _02518_ _02515_ _02519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09178__A2 _04543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07189__A1 _02637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08386__B1 _03969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08925__A2 _04381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05739__A2 _01441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07965_ _03705_ _03693_ _03706_ _00840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09704_ _00098_ io_in[4] u_cpu.rf_ram.memory\[82\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06916_ _03104_ _03100_ _03105_ _00391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07896_ _03500_ _03662_ _03665_ _00812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09635_ _04638_ _04802_ _04810_ _01406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09350__A2 _04641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06847_ _02893_ _03059_ _03065_ _00362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07361__A1 _03312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09566_ u_cpu.rf_ram.memory\[25\]\[0\] _04772_ _04773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06778_ _02897_ _03018_ _03026_ _00332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_70_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10501__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08517_ _04116_ _04117_ _00981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05729_ _02302_ _02304_ u_cpu.cpu.o_wdata1 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09497_ u_cpu.cpu.genblk3.csr.mcause3_0\[2\] _04729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_51_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08861__A1 _03697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07664__A2 _03523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08448_ _04052_ _04056_ _04057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05675__A1 _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08379_ _04000_ _03918_ _03930_ _03944_ _04001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_109_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10410_ _00783_ io_in[4] u_cpu.rf_ram.memory\[91\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10651__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08613__A1 _04013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07416__A2 _03385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05427__A1 _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10341_ _00727_ io_in[4] u_cpu.rf_ram.memory\[125\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05828__I io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09169__A2 _04533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10272_ _00658_ io_in[4] u_cpu.rf_ram.memory\[133\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11007__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08916__A2 _04381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08392__A3 _03962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05450__I1 u_cpu.rf_ram.memory\[49\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10031__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11157__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05038__S0 _01522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09341__A2 _04624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06155__A2 _02637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10181__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05512__B _01519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07655__A2 _03523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05666__A1 _01617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05210__S0 _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10608_ _00981_ io_in[4] u_cpu.cpu.immdec.imm30_25\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07407__A2 _03375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05418__A1 _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08080__A2 _03770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10539_ _00912_ io_in[4] u_cpu.rf_ram.memory\[33\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05738__I _01444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08907__A2 _04371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09580__A2 _04772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06394__A2 _02794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07591__A1 _02632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07750_ u_cpu.rf_ram.memory\[38\]\[4\] _03573_ _03578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04962_ _01543_ _01546_ _01547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09332__A2 _04624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06701_ u_cpu.rf_ram.memory\[129\]\[5\] _02978_ _02984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10524__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07681_ _03506_ _03533_ _03539_ _00722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_04893_ _01474_ _01479_ _01480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07343__A1 _03312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08540__B1 _04004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09420_ _04626_ _04681_ _04683_ _01318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06632_ _02677_ _02695_ _02944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07894__A2 _03662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09351_ u_cpu.rf_ram.memory\[59\]\[3\] _04641_ _04645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06563_ _02666_ _02897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05514_ u_cpu.rf_ram.memory\[4\]\[6\] u_cpu.rf_ram.memory\[5\]\[6\] u_cpu.rf_ram.memory\[6\]\[6\]
+ u_cpu.rf_ram.memory\[7\]\[6\] _01523_ _01525_ _02093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08302_ _03917_ _03919_ _03929_ _03930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_09282_ _04602_ _04603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10674__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06494_ _02685_ _02851_ _02855_ _00219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07646__A2 _03513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08694__I1 u_arbiter.i_wb_cpu_dbus_adr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05657__A1 _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08233_ _02445_ _03874_ _03875_ _00939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05445_ _01543_ _02024_ _02025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05121__A3 _01704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09399__A2 _04671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08164_ _02924_ _03802_ _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05376_ u_cpu.rf_ram.memory\[124\]\[4\] u_cpu.rf_ram.memory\[125\]\[4\] u_cpu.rf_ram.memory\[126\]\[4\]
+ u_cpu.rf_ram.memory\[127\]\[4\] _01496_ _01594_ _01957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__05409__A1 _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07115_ _03098_ _03217_ _03218_ _00477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08095_ _02717_ _02965_ _03779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08071__A2 _03760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06082__A1 _02402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07046_ u_cpu.rf_ram.memory\[58\]\[2\] _03177_ _03180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08359__B1 _03940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09020__A1 _04444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10054__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05268__S0 _01496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09571__A2 _04772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06385__A2 _02784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08997_ _02651_ _04444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07948_ _02636_ _03695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09323__A2 _04624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07879_ u_cpu.rf_ram.memory\[92\]\[3\] _03652_ _03656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09618_ _02619_ _04349_ _04801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07885__A2 _03652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10890_ _01259_ io_in[4] u_cpu.rf_ram.memory\[83\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09549_ _04622_ _04762_ _04763_ _01367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05332__B _01481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07637__A2 _03513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08062__A2 _03760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10324_ _00710_ io_in[4] u_cpu.rf_ram.memory\[127\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10255_ _00641_ io_in[4] u_cpu.rf_ram.memory\[135\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05259__S0 _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09562__A2 _04762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10547__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10186_ _00572_ io_in[4] u_cpu.rf_ram.memory\[71\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06376__A2 _02784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07573__A1 _03306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09314__A2 _04613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07325__A1 _03312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10697__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07876__A2 _03652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07628__A2 _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06300__A2 _02733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07948__I _02636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05230_ u_cpu.rf_ram.memory\[136\]\[2\] u_cpu.rf_ram.memory\[137\]\[2\] u_cpu.rf_ram.memory\[138\]\[2\]
+ u_cpu.rf_ram.memory\[139\]\[2\] _01634_ _01635_ _01813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_144_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05161_ _01737_ _01739_ _01741_ _01743_ _01486_ _01744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__04862__A2 u_cpu.cpu.decode.op26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09250__A1 _04438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08053__A2 _03750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10077__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05498__S0 _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05092_ u_cpu.rf_ram.memory\[60\]\[1\] u_cpu.rf_ram.memory\[61\]\[1\] u_cpu.rf_ram.memory\[62\]\[1\]
+ u_cpu.rf_ram.memory\[63\]\[1\] _01562_ _01563_ _01676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07800__A2 _03605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05811__A1 _02273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08920_ u_cpu.rf_ram.memory\[93\]\[5\] _04381_ _04387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09002__A1 _04446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09553__A2 _04762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08851_ u_cpu.cpu.ctrl.o_ibus_adr\[31\] _04308_ _04329_ _04347_ _04348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_112_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07802_ _02291_ _03605_ _03607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05994_ u_cpu.cpu.ctrl.o_ibus_adr\[12\] _02499_ _02503_ _02504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08782_ _02395_ _02599_ _04310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09305__A2 _04613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07733_ _03504_ _03563_ _03568_ _00745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_04945_ _01529_ _01530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05670__S0 _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08513__B1 _04113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07664_ u_cpu.rf_ram.memory\[127\]\[6\] _03523_ _03530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04876_ _01439_ _01438_ _01462_ _01463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_53_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09403_ u_cpu.rf_ram.memory\[110\]\[2\] _04671_ _04674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06615_ _02934_ _02935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07595_ _02642_ _03485_ _03488_ _00687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_34_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06546_ u_cpu.rf_ram.memory\[50\]\[1\] _02883_ _02886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09334_ _02656_ _04634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07619__A2 _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06477_ _02687_ _02840_ _02845_ _00212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09265_ u_cpu.rf_ram.memory\[83\]\[0\] _04593_ _04594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08216_ u_arbiter.i_wb_cpu_dbus_dat\[20\] _03808_ _03864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05428_ u_cpu.rf_ram.memory\[0\]\[5\] u_cpu.rf_ram.memory\[1\]\[5\] u_cpu.rf_ram.memory\[2\]\[5\]
+ u_cpu.rf_ram.memory\[3\]\[5\] _01530_ _01532_ _02008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09196_ _04438_ _04553_ _04555_ _01222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09712__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08147_ _03810_ _03812_ _02924_ _03813_ _03814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05359_ _01566_ _01939_ _01480_ _01940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_134_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08044__A2 _03750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06055__A1 _02389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05489__S0 _01529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08078_ _03769_ _03770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_49_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07029_ _02642_ _03167_ _03170_ _00439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05802__A1 _02273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08689__I _02335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10040_ _00434_ io_in[4] u_cpu.rf_ram.memory\[19\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09862__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09544__A2 _04752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06358__A2 _02770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07555__A1 _03306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05661__S0 _01507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05046__C _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07307__A1 _03312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10942_ _01311_ io_in[4] u_cpu.rf_ram.memory\[110\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05841__I u_arbiter.i_wb_cpu_dbus_we vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10873_ _01242_ io_in[4] u_cpu.rf_ram.memory\[106\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06530__A2 _02872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09480__A1 _04632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08283__A2 _03910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06294__A1 _02642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09232__A1 _04438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08035__A2 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06046__A1 _02463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06597__A2 _02920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07794__A1 _02263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10307_ _00693_ io_in[4] u_cpu.rf_ram.memory\[22\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09535__A2 _04752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__04920__I _01504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10238_ _00624_ io_in[4] u_cpu.rf_ram.memory\[49\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08594__I0 u_arbiter.i_wb_cpu_rdt\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05237__B _01482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10169_ _00555_ io_in[4] u_cpu.rf_ram.memory\[72\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05652__S0 _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09299__A1 _02675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07849__A2 _03626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06400_ u_cpu.rf_ram.memory\[46\]\[5\] _02794_ _02800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06068__B _02456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07380_ u_cpu.rf_ram.memory\[14\]\[3\] _03365_ _03369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06331_ _02681_ _02756_ _02758_ _00153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09735__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09050_ _02677_ _02814_ _04475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06285__A1 _02728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05088__A2 _01671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06262_ _02693_ _02707_ _02715_ _00127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08001_ u_cpu.rf_ram.memory\[121\]\[6\] _03720_ _03727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05213_ _01597_ _01795_ _01600_ _01796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10712__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08026__A2 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06193_ u_cpu.rf_ram_if.rcnt\[0\] u_cpu.rf_ram_if.rcnt\[1\] _01494_ u_cpu.rf_ram_if.rcnt\[2\]
+ _02670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_116_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05144_ u_cpu.rf_ram.memory\[132\]\[1\] u_cpu.rf_ram.memory\[133\]\[1\] u_cpu.rf_ram.memory\[134\]\[1\]
+ u_cpu.rf_ram.memory\[135\]\[1\] _01634_ _01635_ _01728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09885__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06588__A2 _02912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07785__A1 _03502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09952_ _00346_ io_in[4] u_cpu.rf_ram.memory\[6\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05075_ _01493_ _01658_ _01659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10862__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09526__A2 _03611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08903_ _02657_ _04371_ _04377_ _01107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_106_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09883_ _00277_ io_in[4] u_cpu.rf_ram.memory\[40\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07537__A1 _03306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08834_ u_cpu.cpu.ctrl.o_ibus_adr\[24\] _04327_ _04329_ u_cpu.cpu.ctrl.o_ibus_adr\[25\]
+ _04338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08765_ _03691_ _04299_ _04300_ _01046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05977_ _02403_ u_scanchain_local.module_data_in\[45\] _02478_ u_arbiter.i_wb_cpu_dbus_adr\[8\]
+ _02491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_54_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06760__A2 _03008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07716_ u_cpu.rf_ram.memory\[124\]\[5\] _03553_ _03559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04928_ _01512_ _01513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08696_ u_arbiter.i_wb_cpu_dbus_adr\[5\] u_arbiter.i_wb_cpu_dbus_adr\[6\] _04257_
+ _04261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_65_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07647_ _03508_ _03513_ _03520_ _00707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04859_ _01444_ _01445_ _01446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_53_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06512__A2 _02861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10242__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07578_ u_cpu.rf_ram.memory\[130\]\[3\] _03475_ _03479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09317_ _02631_ _04622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06529_ _02683_ _02872_ _02875_ _00234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09462__A1 _04632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08265__A2 _03885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06276__A1 _02687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05079__A2 _01662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09248_ _04434_ _04583_ _04584_ _01245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10392__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09214__A1 _04438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05874__I1 u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08017__A2 _03730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09179_ u_cpu.rf_ram.memory\[99\]\[2\] _04543_ _04546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06579__A2 _02900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07776__A1 _02717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11141_ _00074_ io_in[0] u_scanchain_local.module_data_in\[53\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05836__I _02395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05251__A2 _01832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11072_ _01432_ io_in[4] u_cpu.rf_ram_if.rdata1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10023_ _00417_ io_in[4] u_cpu.rf_ram.memory\[61\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06751__A2 _03008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10925_ _01294_ io_in[4] u_cpu.rf_ram.memory\[10\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09758__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06503__A2 _02827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10856_ _01225_ io_in[4] u_cpu.rf_ram.memory\[79\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10735__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08256__A2 _03885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10787_ _01156_ io_in[4] u_cpu.cpu.genblk1.align.ctrl_misal vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__04915__I _01499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08008__A2 _03730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06019__A1 _02388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10885__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05490__A2 _02069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07767__A1 _03502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05242__A2 _01823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10115__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07519__A1 _03306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06990__A2 _03147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05900_ _02436_ _00041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06880_ u_cpu.rf_ram.memory\[65\]\[4\] _03079_ _03084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05831_ _01441_ _02355_ _02260_ _02306_ _02391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_67_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08319__I0 u_arbiter.i_wb_cpu_rdt\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06742__A2 _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10265__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08550_ _04141_ _04142_ _04147_ _00984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05762_ _02322_ _02323_ _02337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07501_ _03306_ _03435_ _03436_ _00645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05693_ _02263_ u_cpu.cpu.immdec.imm31 _02269_ _02270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08481_ _04069_ _04083_ _04084_ _04085_ _00977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__05414__C _01466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08495__A2 _04097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09692__A1 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07432_ u_cpu.rf_ram.memory\[137\]\[2\] _03395_ _03398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08247__A2 _03835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07363_ _03314_ _03355_ _03359_ _00584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09444__A1 _04632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09102_ _04502_ _04503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06258__A1 _02689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06314_ _02642_ _02745_ _02748_ _00146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07294_ _02661_ _03320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09033_ u_cpu.rf_ram.memory\[96\]\[2\] _04463_ _04466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06245_ _02619_ _02677_ _02706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05481__A2 _02060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06176_ _02655_ _02656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07758__A1 _02675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05127_ _01602_ _01710_ _01711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05233__A2 _01815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09935_ _00329_ io_in[4] u_cpu.rf_ram.memory\[76\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05058_ u_cpu.rf_ram.memory\[128\]\[0\] u_cpu.rf_ram.memory\[129\]\[0\] u_cpu.rf_ram.memory\[130\]\[0\]
+ u_cpu.rf_ram.memory\[131\]\[0\] _01641_ _01642_ _01643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__11040__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06981__A2 _03137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09866_ _00260_ io_in[4] u_cpu.raddr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10608__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08817_ _04310_ _04329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09797_ _00191_ io_in[4] u_cpu.rf_ram.memory\[45\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06733__A2 _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07930__A1 _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09900__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05092__S1 _01563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08748_ _02590_ _02592_ _02598_ _04287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05605__B _01534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10758__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09683__A1 _04632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08679_ u_cpu.rf_ram.memory\[31\]\[4\] _04247_ _04252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08486__A2 _03940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10710_ _01080_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10641_ _01014_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10572_ _00945_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10138__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07749__A1 _03502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08410__A2 _04020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05224__A2 _01806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11124_ _00055_ io_in[0] u_scanchain_local.module_data_in\[36\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06972__A2 _03137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10288__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11055_ _01423_ io_in[4] u_cpu.rf_ram.memory\[23\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08174__A1 u_arbiter.i_wb_cpu_dbus_dat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10006_ _00400_ io_in[4] u_cpu.rf_ram.memory\[63\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06724__A2 _02988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05083__S1 _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06488__A1 _02669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10908_ _01277_ io_in[4] u_cpu.rf_ram.memory\[84\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09426__A1 _04632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10839_ _01208_ io_in[4] u_cpu.rf_ram.memory\[104\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05160__A1 _01506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08229__A2 _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06030_ u_arbiter.i_wb_cpu_dbus_adr\[19\] _02397_ _02533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05463__A2 _02038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06660__A1 _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11063__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05215__A2 _01797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06412__A1 _02681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07981_ u_cpu.rf_ram.memory\[118\]\[5\] _03710_ _03716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08952__A3 _02604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06963__A2 _03127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09720_ _00114_ io_in[4] u_cpu.rf_ram.memory\[81\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09923__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06932_ _02827_ _02870_ _03116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__04974__A1 _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09651_ _04636_ _04812_ _04819_ _01413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06863_ _02891_ _03069_ _03074_ _00369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10900__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06715__A2 _02988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07912__A1 _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08602_ _03928_ _03986_ _04177_ _04193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__05074__S1 _01525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05814_ u_cpu.rf_ram_if.rdata0\[1\] _01467_ _02381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09582_ _02677_ _02954_ _04781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06794_ _02895_ _03028_ _03035_ _00339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08533_ _03908_ _04131_ _04079_ _03910_ _04132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_36_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05745_ u_cpu.cpu.immdec.imm31 _02269_ _02320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09665__A1 _04632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08468__A2 _04068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06479__A1 _02689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08464_ _04019_ _04071_ _00974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05676_ u_cpu.rf_ram.memory\[136\]\[7\] u_cpu.rf_ram.memory\[137\]\[7\] u_cpu.rf_ram.memory\[138\]\[7\]
+ u_cpu.rf_ram.memory\[139\]\[7\] _01641_ _01642_ _02254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07140__A2 _03227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07415_ _03312_ _03385_ _03388_ _00607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05151__A1 _01725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08395_ _03899_ _03988_ _04015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05160__B _01519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07346_ u_cpu.rf_ram.memory\[70\]\[4\] _03345_ _03350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07277_ u_cpu.rf_ram.memory\[72\]\[0\] _03308_ _03309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08640__A2 _02320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09016_ _04440_ _04453_ _04456_ _01141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06651__A1 _02782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05454__A2 _02005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06228_ _02696_ _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06159_ _02641_ _02642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10430__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06403__A1 _02691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08943__A3 _03985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06954__A2 _03127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09918_ _00312_ io_in[4] u_cpu.rf_ram.memory\[77\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__04965__A1 _01548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09849_ _00243_ io_in[4] u_cpu.rf_ram.memory\[50\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10580__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06706__A2 _02978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05065__S1 _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08459__A2 _03956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09408__A1 _04632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10624_ _00997_ io_in[4] u_cpu.rf_ram.memory\[32\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05693__A2 u_cpu.cpu.immdec.imm31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11086__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10555_ _00928_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08631__A2 _04165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05445__A2 _02024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10486_ _00859_ io_in[4] u_cpu.rf_ram.memory\[8\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09946__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08395__A1 _03899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07198__A2 _03257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06945__A2 _03117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10923__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11107_ _00036_ io_in[0] u_arbiter.i_wb_cpu_rdt\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05599__I3 u_cpu.rf_ram.memory\[19\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11038_ _01407_ io_in[4] u_cpu.rf_ram.memory\[100\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07370__A2 _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09647__A1 _04632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05381__A1 _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05530_ _01463_ _02108_ _01558_ _02109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_75_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07122__A2 _03217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10303__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05461_ u_cpu.rf_ram.memory\[104\]\[5\] u_cpu.rf_ram.memory\[105\]\[5\] u_cpu.rf_ram.memory\[106\]\[5\]
+ u_cpu.rf_ram.memory\[107\]\[5\] _01555_ _01531_ _02041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_32_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08870__A2 _04351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07200_ u_cpu.rf_ram.memory\[15\]\[7\] _03257_ _03265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05684__A2 u_cpu.cpu.bufreg.i_sh_signed vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06881__A1 _02891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05392_ u_cpu.rf_ram.memory\[84\]\[4\] u_cpu.rf_ram.memory\[85\]\[4\] u_cpu.rf_ram.memory\[86\]\[4\]
+ u_cpu.rf_ram.memory\[87\]\[4\] _01507_ _01605_ _01973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08180_ u_arbiter.i_wb_cpu_dbus_dat\[8\] _03835_ _03840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07131_ _03226_ _03227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10453__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05436__A2 _02015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07062_ u_cpu.rf_ram.memory\[57\]\[1\] _03187_ _03189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06013_ u_cpu.cpu.ctrl.o_ibus_adr\[16\] _02518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_12_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08386__A1 _03974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07189__A2 _03257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05139__C _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06936__A2 _03117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07964_ u_cpu.rf_ram.memory\[120\]\[6\] _03693_ _03706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09703_ _00097_ io_in[4] u_cpu.rf_ram.memory\[82\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06915_ u_cpu.rf_ram.memory\[29\]\[2\] _03100_ _03105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07895_ u_cpu.rf_ram.memory\[35\]\[2\] _03662_ _03665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09634_ u_cpu.rf_ram.memory\[98\]\[7\] _04802_ _04810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06846_ u_cpu.rf_ram.memory\[67\]\[5\] _03059_ _03065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05870__S _02418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07361__A2 _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05372__A1 _01512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09565_ _04771_ _04772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06777_ u_cpu.rf_ram.memory\[76\]\[7\] _03018_ _03026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08516_ u_cpu.cpu.immdec.imm30_25\[2\] _04104_ _04106_ u_cpu.cpu.immdec.imm30_25\[3\]
+ _04113_ _04009_ _04117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_05728_ u_arbiter.i_wb_cpu_ibus_adr\[0\] _02303_ _02304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09819__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09496_ _02295_ _04723_ _04728_ _01349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08310__A1 _02466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08447_ _04024_ _04054_ _04055_ _04056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05659_ u_cpu.rf_ram.memory\[64\]\[7\] u_cpu.rf_ram.memory\[65\]\[7\] u_cpu.rf_ram.memory\[66\]\[7\]
+ u_cpu.rf_ram.memory\[67\]\[7\] _01522_ _01622_ _02237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08861__A2 _04351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05675__A2 _02252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08378_ u_arbiter.i_wb_cpu_rdt\[12\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[12\]
+ _02466_ _04000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09969__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07329_ _03316_ _03335_ _03340_ _00569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08613__A2 _04052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10340_ _00726_ io_in[4] u_cpu.rf_ram.memory\[125\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10946__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10271_ _00657_ io_in[4] u_cpu.rf_ram.memory\[133\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06927__A2 _03100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05844__I _02402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05038__S1 _01622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07352__A2 _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10326__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09629__A1 _04632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05363__A1 _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07104__A2 _03207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05115__A1 _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10476__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05210__S1 _01563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05666__A2 _02243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06863__A1 _02891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10607_ _00980_ io_in[4] u_cpu.cpu.immdec.imm30_25\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05418__A2 _01997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04923__I _01507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10538_ _00911_ io_in[4] u_cpu.rf_ram.memory\[33\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10469_ _00842_ io_in[4] u_cpu.rf_ram.memory\[118\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08368__A1 _03915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06918__A2 _03100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07040__A1 _02780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11101__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07591__A2 _03485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04961_ u_cpu.rf_ram.memory\[36\]\[0\] u_cpu.rf_ram.memory\[37\]\[0\] u_cpu.rf_ram.memory\[38\]\[0\]
+ u_cpu.rf_ram.memory\[39\]\[0\] _01544_ _01545_ _01546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_06700_ _02891_ _02978_ _02983_ _00297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07680_ u_cpu.rf_ram.memory\[126\]\[5\] _03533_ _03539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04892_ _01475_ _01452_ _01476_ _01447_ _01478_ _01479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_64_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08540__A1 _03922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07343__A2 _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06631_ _02897_ _02935_ _02943_ _00268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_93_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05354__A1 _01463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09350_ _04628_ _04641_ _04644_ _01287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10819__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06562_ _02895_ _02883_ _02896_ _00246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08301_ _03926_ _03928_ _03929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05513_ _02085_ _02087_ _02089_ _02091_ _01486_ _02092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__05106__A1 _01548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09281_ _02814_ _04349_ _04602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06493_ u_cpu.rf_ram.memory\[43\]\[3\] _02851_ _02855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05657__A2 _02234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08232_ u_arbiter.i_wb_cpu_rdt\[25\] _03807_ _03808_ u_arbiter.i_wb_cpu_dbus_dat\[25\]
+ _03875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05444_ u_cpu.rf_ram.memory\[60\]\[5\] u_cpu.rf_ram.memory\[61\]\[5\] u_cpu.rf_ram.memory\[62\]\[5\]
+ u_cpu.rf_ram.memory\[63\]\[5\] _01496_ _01594_ _02024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_119_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05901__I0 u_arbiter.i_wb_cpu_rdt\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10969__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08163_ _02915_ _03826_ _03827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05375_ _01949_ _01951_ _01953_ _01955_ _01560_ _01956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__05409__A2 _01989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07114_ u_cpu.rf_ram.memory\[54\]\[0\] _03217_ _03218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08094_ _03707_ _03770_ _03778_ _00897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07045_ _03102_ _03177_ _03179_ _00446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_47_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08359__A1 _02305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08359__B2 _03959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09020__A2 _04453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06909__A2 _03100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07031__A1 _02647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05268__S1 _01563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08996_ _04442_ _04436_ _04443_ _01134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07582__A2 _03475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10349__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07947_ _03691_ _03693_ _03694_ _00834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07878_ _03500_ _03652_ _03655_ _00804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_18_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07334__A2 _03335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09617_ _02693_ _04792_ _04800_ _01398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_83_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05345__A1 _01513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06829_ _02893_ _03049_ _03055_ _00354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10499__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09548_ u_cpu.rf_ram.memory\[26\]\[0\] _04762_ _04763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09479_ u_cpu.rf_ram.memory\[88\]\[4\] _04711_ _04716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09791__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08834__A2 _04327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05648__A2 _02221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06845__A1 _02891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__04951__S0 _01523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08598__A1 _03940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10323_ _00709_ io_in[4] u_cpu.rf_ram.memory\[127\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06073__A2 _02562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11124__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10254_ _00640_ io_in[4] u_cpu.rf_ram.memory\[135\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05820__A2 _01467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09011__A2 _04453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07022__A1 _02675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05259__S1 _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10185_ _00571_ io_in[4] u_cpu.rf_ram.memory\[71\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07573__A2 _03475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08522__A1 _03924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06128__A3 _02612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07325__A2 _03335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05336__A1 _01506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07089__A1 _03110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05639__A2 _02212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05195__S0 _01529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05160_ _01506_ _01742_ _01519_ _01743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09250__A2 _04583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07261__A1 _02637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05498__S1 _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05091_ _01668_ _01670_ _01672_ _01674_ _01560_ _01675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_144_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09002__A2 _04436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07013__A1 _03106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08850_ _01451_ _04345_ _04346_ _04347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_112_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07801_ _02291_ _03605_ _03606_ _00775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07564__A2 _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08781_ _04308_ _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05993_ u_cpu.cpu.ctrl.o_ibus_adr\[12\] _02499_ _02461_ _02503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07732_ u_cpu.rf_ram.memory\[123\]\[4\] _03563_ _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04944_ _01494_ _01529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__05670__S1 _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10641__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08513__A1 _03932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07316__A2 _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08513__B2 _03909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07663_ _03506_ _03523_ _03529_ _00714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05327__A1 _01899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04875_ _01453_ _01461_ _01462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_65_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07867__A3 _02291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09402_ _04626_ _04671_ _04673_ _01310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06614_ _02677_ _02754_ _02934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05433__B _01482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07594_ u_cpu.rf_ram.memory\[12\]\[2\] _03485_ _03488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09333_ _04632_ _04624_ _04633_ _01281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10791__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06545_ _02636_ _02885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06827__A1 _02891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09264_ _04592_ _04593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06476_ u_cpu.rf_ram.memory\[41\]\[4\] _02840_ _02845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05186__S0 _01576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08215_ _03862_ _03863_ _00933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05427_ _01493_ _02006_ _02007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09195_ u_cpu.rf_ram.memory\[79\]\[1\] _04553_ _04555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10021__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11147__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08146_ u_arbiter.i_wb_cpu_dbus_dat\[1\] _03804_ _03813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05358_ u_cpu.rf_ram.memory\[56\]\[4\] u_cpu.rf_ram.memory\[57\]\[4\] u_cpu.rf_ram.memory\[58\]\[4\]
+ u_cpu.rf_ram.memory\[59\]\[4\] _01567_ _01568_ _01939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09241__A2 _04573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08077_ _02825_ _02965_ _03769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05489__S1 _01500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05289_ _01543_ _01870_ _01871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07028_ u_cpu.rf_ram.memory\[5\]\[2\] _03167_ _03170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_1_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10171__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07004__A1 _02677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07555__A2 _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08979_ u_cpu.rf_ram.memory\[97\]\[6\] _04425_ _04432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05661__S1 _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08504__A1 _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07307__A2 _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10941_ _01310_ io_in[4] u_cpu.rf_ram.memory\[110\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10872_ _01241_ io_in[4] u_cpu.rf_ram.memory\[106\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05062__C _01466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05177__S0 _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09480__A2 _04711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07491__A1 _03316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06294__A2 _02733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09232__A2 _04573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10514__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07243__A1 _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07794__A2 _02914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10306_ _00692_ io_in[4] u_cpu.rf_ram.memory\[12\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10237_ _00623_ io_in[4] u_cpu.rf_ram.memory\[49\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10664__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07546__A2 _03455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08594__I1 u_arbiter.i_wb_cpu_rdt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05557__A1 _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10168_ _00554_ io_in[4] u_cpu.rf_ram.memory\[72\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05652__S1 _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10099_ _00493_ io_in[4] u_cpu.rf_ram.memory\[52\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09299__A2 _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08548__C _02585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05253__B _01534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10044__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08564__B _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06809__A1 _02652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06330_ u_cpu.rf_ram.memory\[80\]\[1\] _02756_ _02758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05168__S0 _01530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09471__A2 _04711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06285__A2 _02608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06261_ u_cpu.rf_ram.memory\[18\]\[7\] _02707_ _02715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08000_ _03703_ _03720_ _03726_ _00855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05212_ u_cpu.rf_ram.memory\[88\]\[2\] u_cpu.rf_ram.memory\[89\]\[2\] u_cpu.rf_ram.memory\[90\]\[2\]
+ u_cpu.rf_ram.memory\[91\]\[2\] _01598_ _01556_ _01795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_11_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06192_ _02631_ _02669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10194__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09223__A2 _04563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05143_ _01465_ _01726_ _01727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08982__A1 _03707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07785__A2 _03593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05074_ u_cpu.rf_ram.memory\[4\]\[1\] u_cpu.rf_ram.memory\[5\]\[1\] u_cpu.rf_ram.memory\[6\]\[1\]
+ u_cpu.rf_ram.memory\[7\]\[1\] _01523_ _01525_ _01658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09951_ _00345_ io_in[4] u_cpu.rf_ram.memory\[6\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05796__A1 _02273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05340__S0 _01530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08902_ u_cpu.rf_ram.memory\[2\]\[5\] _04371_ _04377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09882_ _00276_ io_in[4] u_cpu.rf_ram.memory\[17\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07537__A2 _03455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08833_ _04337_ _01077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05548__A1 _01512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08764_ u_cpu.rf_ram.memory\[30\]\[0\] _04299_ _04300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05976_ _02456_ _02489_ _02490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07715_ _03504_ _03553_ _03558_ _00737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04927_ _01463_ _01512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_54_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08695_ _04260_ _01016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07646_ u_cpu.rf_ram.memory\[128\]\[6\] _03513_ _03520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04858_ u_cpu.cpu.branch_op _01445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_81_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05720__A1 _02263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07577_ _03312_ _03475_ _03478_ _00679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09316_ _04450_ _04613_ _04621_ _01276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06528_ u_cpu.rf_ram.memory\[47\]\[2\] _02872_ _02875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05159__S0 _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09462__A2 _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10537__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09247_ u_cpu.rf_ram.memory\[107\]\[0\] _04583_ _04584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06276__A2 _02719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07473__A1 _03316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05610__C _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06459_ u_cpu.rf_ram.memory\[51\]\[5\] _02829_ _02835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09178_ _04438_ _04543_ _04545_ _01214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09214__A2 _04563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07225__A1 _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08129_ u_cpu.rf_ram.memory\[33\]\[7\] _03790_ _03798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10687__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07776__A2 _02782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11140_ _00073_ io_in[0] u_scanchain_local.module_data_in\[52\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05331__S0 _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11071_ u_cpu.rf_ram_if.wtrig0 io_in[4] u_cpu.rf_ram_if.genblk1.wtrig0_r vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07528__A2 _03445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10022_ _00416_ io_in[4] u_cpu.rf_ram.memory\[61\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05539__A1 _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10067__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09150__A1 _04446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10924_ _01293_ io_in[4] u_cpu.rf_ram.memory\[10\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07700__A2 _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10855_ _01224_ io_in[4] u_cpu.rf_ram.memory\[79\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05711__A1 _02285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10786_ _01155_ io_in[4] u_cpu.cpu.bufreg.i_sh_signed vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09453__A2 _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06267__A2 _02719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09205__A2 _04553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05227__B1 _01807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08964__A1 _02621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07767__A2 _03583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05322__S0 _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05248__B _01519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07519__A2 _03445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08192__A2 _03835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05830_ io_in[2] _02389_ _02390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08319__I1 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05761_ _02306_ _02335_ _02336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09702__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07500_ u_cpu.rf_ram.memory\[134\]\[0\] _03435_ _03436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08480_ u_cpu.cpu.immdec.imm24_20\[3\] _04069_ _04085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05692_ _01444_ _01445_ _01442_ _02269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_74_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07431_ _03310_ _03395_ _03397_ _00614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05702__A1 u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07362_ u_cpu.rf_ram.memory\[143\]\[3\] _03355_ _03359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09852__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09444__A2 _04691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09101_ _02675_ _04349_ _04502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06313_ u_cpu.rf_ram.memory\[7\]\[2\] _02745_ _02748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06258__A2 _02707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07455__A1 _03316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07293_ _03318_ _03308_ _03319_ _00554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09032_ _04438_ _04463_ _04465_ _01148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06244_ _02693_ _02697_ _02705_ _00119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07207__A1 _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06175_ _02611_ u_cpu.rf_ram_if.wdata0_r\[5\] _02654_ _02655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_144_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07758__A2 _02782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05126_ u_cpu.rf_ram.memory\[80\]\[1\] u_cpu.rf_ram.memory\[81\]\[1\] u_cpu.rf_ram.memory\[82\]\[1\]
+ u_cpu.rf_ram.memory\[83\]\[1\] _01496_ _01594_ _01710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_85_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05313__S0 _01529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05769__A1 u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09934_ _00328_ io_in[4] u_cpu.rf_ram.memory\[76\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06430__A2 _02816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05057_ _01622_ _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09865_ _00259_ io_in[4] u_cpu.raddr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08183__A2 _03835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08816_ _04328_ _01069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_09796_ _00190_ io_in[4] u_cpu.rf_ram.memory\[45\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06194__A1 _01498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07930__A2 _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08747_ _04286_ _01042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05959_ _02464_ u_cpu.cpu.ctrl.o_ibus_adr\[4\] u_cpu.cpu.ctrl.o_ibus_adr\[3\] u_cpu.cpu.ctrl.o_ibus_adr\[2\]
+ _02476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_38_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09132__A1 _04446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08983__I _02631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08678_ _03699_ _04247_ _04251_ _01008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09683__A2 _04832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07629_ _02666_ _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06497__A2 _02851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10640_ _01013_ io_in[4] u_cpu.cpu.alu.cmp_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09435__A2 _04691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07446__A1 u_cpu.rf_ram.memory\[49\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06249__A2 _02707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10571_ _00944_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07997__A2 _03720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05552__S0 _01496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08946__A1 _03940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07749__A2 _03573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05304__S0 _01507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11123_ _00054_ io_in[0] u_scanchain_local.module_data_in\[35\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05068__B _01481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06421__A2 _02805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11054_ _00025_ io_in[4] u_cpu.rf_ram.regzero vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09725__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08174__A2 _03835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10005_ _00399_ io_in[4] u_cpu.rf_ram.memory\[63\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06185__A1 _02628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07921__A2 _03672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10702__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05932__A1 _02403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09875__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09674__A2 _04832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06488__A2 _02851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07685__A1 _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10907_ _01276_ io_in[4] u_cpu.rf_ram.memory\[69\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10838_ _01207_ io_in[4] u_cpu.rf_ram.memory\[104\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10852__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05160__A2 _01742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09426__A2 _04681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07437__A1 _03316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10769_ _01138_ io_in[4] u_cpu.rf_ram.memory\[94\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05543__S0 _01551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06660__A2 _02956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08937__A1 u_cpu.cpu.immdec.imm11_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06412__A2 _02805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07980_ _03701_ _03710_ _03715_ _00846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10232__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06931_ _03114_ _03100_ _03115_ _00396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09650_ u_cpu.rf_ram.memory\[100\]\[6\] _04812_ _04819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06862_ u_cpu.rf_ram.memory\[66\]\[4\] _03069_ _03074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08601_ _03928_ _04188_ _04189_ _04191_ _03969_ _04192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_110_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05813_ _02272_ _02379_ _02380_ _00020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07912__A2 _03672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09581_ _04638_ _04772_ _04780_ _01382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10382__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05425__C _01486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06793_ u_cpu.rf_ram.memory\[75\]\[6\] _03028_ _03035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09114__A1 _04446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08532_ u_arbiter.i_wb_cpu_rdt\[29\] u_arbiter.i_wb_cpu_rdt\[13\] _02467_ _04131_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05744_ _01445_ _02318_ _02319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_70_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09665__A2 _04822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08712__I1 u_arbiter.i_wb_cpu_dbus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08463_ u_cpu.cpu.immdec.imm24_20\[0\] _04069_ _04070_ u_cpu.cpu.immdec.imm24_20\[1\]
+ _04071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06479__A2 _02840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05675_ _01638_ _02252_ _02253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_35_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07414_ u_cpu.rf_ram.memory\[39\]\[2\] _03385_ _03388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08394_ _03901_ _04012_ _04013_ _04014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_50_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09417__A2 _04681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05151__A2 _01734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07345_ _03314_ _03345_ _03349_ _00576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07979__A2 _03710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05868__S _02418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06100__A1 _02322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07276_ _03307_ _03308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05534__S0 _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09015_ u_cpu.rf_ram.memory\[95\]\[2\] _04453_ _04456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06227_ _02626_ _02695_ _02696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06651__A2 _02954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05454__A3 _02014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08928__A1 u_cpu.cpu.immdec.imm11_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06158_ _02640_ _02641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09748__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05109_ u_cpu.rf_ram.memory\[104\]\[1\] u_cpu.rf_ram.memory\[105\]\[1\] u_cpu.rf_ram.memory\[106\]\[1\]
+ u_cpu.rf_ram.memory\[107\]\[1\] _01555_ _01531_ _01693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06403__A2 _02794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06089_ u_arbiter.i_wb_cpu_dbus_adr\[30\] _02397_ _02578_ _02580_ _02402_ _02581_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_137_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09075__S _04485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09917_ _00311_ io_in[4] u_cpu.rf_ram.memory\[77\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04965__A2 _01549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10725__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09848_ _00242_ io_in[4] u_cpu.rf_ram.memory\[50\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06167__A1 _02628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09898__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07903__A2 _03662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09779_ _00173_ io_in[4] u_cpu.rf_ram.memory\[42\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10875__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09656__A2 _04822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07667__A1 _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09408__A2 _04671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10105__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10623_ _00996_ io_in[4] u_cpu.cpu.genblk3.csr.timer_irq_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07419__A1 _03316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06890__A2 _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08092__A1 _03705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10554_ _00927_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05525__S0 _01495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08381__C _03955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06642__A2 _02945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10485_ _00858_ io_in[4] u_cpu.rf_ram.memory\[8\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10255__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08919__A1 _03701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08395__A2 _03988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11106_ _00035_ io_in[0] u_arbiter.i_wb_cpu_rdt\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11037_ _01406_ io_in[4] u_cpu.rf_ram.memory\[98\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05526__B _01518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09647__A2 _04812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05381__A2 _01961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05460_ _01512_ _02039_ _02040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11030__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05391_ _01602_ _01971_ _01972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06881__A2 _03079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07130_ _02675_ _02827_ _03226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05516__S0 _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07061_ _03098_ _03187_ _03188_ _00453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07830__A1 _03508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06012_ _02456_ _02516_ _02517_ _00075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_126_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10748__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08386__A2 _03904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06397__A1 _02685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07963_ _02661_ _03705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08138__A2 _02397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09702_ _00096_ io_in[4] u_cpu.rf_ram.memory\[82\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06914_ _02641_ _03104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10898__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06149__A1 _02628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07894_ _03498_ _03662_ _03664_ _00811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09633_ _04636_ _04802_ _04809_ _01405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06845_ _02891_ _03059_ _03064_ _00361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09564_ _02677_ _02838_ _04771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06776_ _02895_ _03018_ _03025_ _00331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05372__A2 _01952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09638__A2 _04812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10128__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08515_ _04110_ _04115_ _04116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05727_ u_cpu.cpu.state.genblk1.misalign_trap_sync_r _01459_ _02303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__07649__A1 _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08846__B1 _04329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09495_ _04723_ _04727_ _04728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_24_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08446_ _03922_ _03996_ _04000_ _03998_ _04055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_05658_ _02229_ _02231_ _02233_ _02235_ _01581_ _02236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_51_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06872__A2 _03079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08377_ _03996_ _03940_ _03998_ _03922_ _03999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_104_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05589_ _01638_ _02167_ _01534_ _02168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10278__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04883__A1 u_cpu.cpu.immdec.imm24_20\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07328_ u_cpu.rf_ram.memory\[71\]\[4\] _03335_ _03340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08074__A1 _03705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05507__S0 _01522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06624__A2 _02935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07259_ _02632_ _03297_ _03298_ _00541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10270_ _00656_ io_in[4] u_cpu.rf_ram.memory\[133\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08702__S _04257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08377__A2 _03940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06388__A1 _02766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08129__A2 _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07888__A1 _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09629__A2 _04802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11053__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08301__A2 _03928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05081__B _01482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05115__A2 _01698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06312__A1 _02637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09913__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06863__A2 _03069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10606_ _00979_ io_in[4] u_cpu.cpu.immdec.imm30_25\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07812__A1 _02395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10537_ _00910_ io_in[4] u_cpu.rf_ram.memory\[33\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10468_ _00841_ io_in[4] u_cpu.rf_ram.memory\[120\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06379__A1 _02685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10399_ _00772_ io_in[4] u_cpu.rf_ram.memory\[36\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07040__A2 _02827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04960_ _01499_ _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04891_ _01438_ _01477_ _01478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_49_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06000__B1 _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08540__A2 _03923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06630_ u_cpu.rf_ram.memory\[16\]\[7\] _02935_ _02943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06561_ u_cpu.rf_ram.memory\[50\]\[6\] _02883_ _02896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08828__B1 _04329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08300_ _02909_ u_arbiter.i_wb_cpu_rdt\[8\] _03927_ _03928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_61_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05512_ _01506_ _02090_ _01519_ _02091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10420__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09280_ _04450_ _04593_ _04601_ _01260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06492_ _02683_ _02851_ _02854_ _00218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08231_ _02924_ _03802_ _03874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05443_ _02016_ _02018_ _02020_ _02022_ _01560_ _02023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__06854__A2 _03069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08056__A1 _03705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08162_ u_arbiter.i_wb_cpu_dbus_dat\[4\] _02916_ _03826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05374_ _01566_ _01954_ _01558_ _01955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10570__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07113_ _03216_ _03217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08093_ u_cpu.rf_ram.memory\[115\]\[7\] _03770_ _03778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07803__A1 u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07044_ u_cpu.rf_ram.memory\[58\]\[1\] _03177_ _03179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08359__A2 _03956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05945__I _02464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07031__A2 _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08995_ u_cpu.rf_ram.memory\[94\]\[3\] _04436_ _04443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09308__A1 _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07946_ u_cpu.rf_ram.memory\[120\]\[0\] _03693_ _03694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06790__A1 _02891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08516__C1 _04113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11076__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07877_ u_cpu.rf_ram.memory\[92\]\[2\] _03652_ _03655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09616_ u_cpu.rf_ram.memory\[0\]\[7\] _04792_ _04800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_16_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06828_ u_cpu.rf_ram.memory\[68\]\[5\] _03049_ _03055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09547_ _04761_ _04762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06759_ u_cpu.rf_ram.memory\[74\]\[7\] _03008_ _03016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09936__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07098__A2 _03207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08991__I _02641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09478_ _04630_ _04711_ _04715_ _01344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_93_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08429_ u_cpu.rf_ram.memory\[114\]\[2\] _04041_ _04044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06845__A2 _03059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10913__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__04856__A1 _01441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09095__I0 u_arbiter.i_wb_cpu_rdt\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04951__S1 _01525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08598__A2 _03929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10322_ _00708_ io_in[4] u_cpu.rf_ram.memory\[128\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07270__A2 _03297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10253_ _00639_ io_in[4] u_cpu.rf_ram.memory\[135\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07022__A2 _02731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10184_ _00570_ io_in[4] u_cpu.rf_ram.memory\[71\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08770__A2 _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08522__A2 _03910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10443__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05336__A2 _01916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06533__A1 _02687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08286__A1 _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07089__A2 _03197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10593__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06836__A2 _03059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05195__S1 _01524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05895__I0 u_arbiter.i_wb_cpu_rdt\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08038__A1 _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04934__I _01518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05090_ _01554_ _01673_ _01558_ _01674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07261__A2 _03297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09809__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07013__A2 _03157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11099__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07800_ _02291_ _03605_ _02396_ _03606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08780_ _02259_ _02598_ _02395_ _04308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_57_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05992_ _02502_ _00069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_69_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06772__A1 _02891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07731_ _03502_ _03563_ _03567_ _00744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_04943_ _01505_ _01528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_66_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09959__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08513__A2 _04051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07662_ u_cpu.rf_ram.memory\[127\]\[5\] _03523_ _03529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04874_ _01455_ _01456_ u_cpu.rf_ram_if.rtrig0 _01460_ _01461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_66_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05327__A2 _01908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09401_ u_cpu.rf_ram.memory\[110\]\[1\] _04671_ _04673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06613_ _02928_ _02933_ _00260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_77_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07593_ _02637_ _03485_ _03487_ _00686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10936__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09332_ u_cpu.rf_ram.memory\[84\]\[4\] _04624_ _04633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06544_ _02881_ _02883_ _02884_ _00240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09263_ _02626_ _02825_ _04592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06475_ _02685_ _02840_ _02844_ _00211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06827__A2 _03049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05186__S1 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08214_ u_arbiter.i_wb_cpu_rdt\[19\] _03807_ _03829_ u_arbiter.i_wb_cpu_dbus_dat\[20\]
+ _03863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__05886__I0 u_arbiter.i_wb_cpu_rdt\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05426_ u_cpu.rf_ram.memory\[4\]\[5\] u_cpu.rf_ram.memory\[5\]\[5\] u_cpu.rf_ram.memory\[6\]\[5\]
+ u_cpu.rf_ram.memory\[7\]\[5\] _01523_ _01525_ _02006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_119_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09194_ _04434_ _04553_ _04554_ _01221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09077__I0 u_arbiter.i_wb_cpu_rdt\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08145_ _03802_ _03811_ _03812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05357_ _01464_ _01937_ _01938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05876__S _02418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08076_ _03707_ _03760_ _03768_ _00889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07252__A2 _03287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05288_ u_cpu.rf_ram.memory\[124\]\[3\] u_cpu.rf_ram.memory\[125\]\[3\] u_cpu.rf_ram.memory\[126\]\[3\]
+ u_cpu.rf_ram.memory\[127\]\[3\] _01496_ _01594_ _01870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10316__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07027_ _02637_ _03167_ _03169_ _00438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_115_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07004__A2 _02825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10466__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08978_ _03703_ _04425_ _04431_ _01128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09083__S _04485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07929_ u_cpu.rf_ram.memory\[117\]\[1\] _03682_ _03684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08504__A2 _04101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09701__A1 _02927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10940_ _01309_ io_in[4] u_cpu.rf_ram.memory\[110\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10871_ _01240_ io_in[4] u_cpu.rf_ram.memory\[106\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06818__A2 _03049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05177__S1 _01531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07491__A2 _03425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08440__A1 _03707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07243__A2 _03287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10305_ _00691_ io_in[4] u_cpu.rf_ram.memory\[12\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10809__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10236_ _00622_ io_in[4] u_cpu.rf_ram.memory\[49\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10167_ _00553_ io_in[4] u_cpu.rf_ram.memory\[72\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05557__A2 _02135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06754__A1 _02891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10098_ _00492_ io_in[4] u_cpu.rf_ram.memory\[53\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10959__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06506__A1 _02669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08259__A1 _03701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06809__A2 _03039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05168__S1 _01532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05868__I0 u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06260_ _02691_ _02707_ _02714_ _00126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07482__A2 _03425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10339__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05211_ _01464_ _01793_ _01794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05493__A1 _02053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06191_ _02628_ _02667_ _02668_ _00103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05142_ u_cpu.rf_ram.memory\[128\]\[1\] u_cpu.rf_ram.memory\[129\]\[1\] u_cpu.rf_ram.memory\[130\]\[1\]
+ u_cpu.rf_ram.memory\[131\]\[1\] _01634_ _01635_ _01726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07234__A2 _03277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08982__A2 _04425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05073_ _01650_ _01652_ _01654_ _01656_ _01486_ _01657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_09950_ _00344_ io_in[4] u_cpu.rf_ram.memory\[6\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10489__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06993__A1 _03104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05340__S1 _01532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08901_ _02652_ _04371_ _04376_ _01106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_98_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09881_ _00275_ io_in[4] u_cpu.rf_ram.memory\[17\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09781__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08832_ u_cpu.cpu.ctrl.o_ibus_adr\[23\] _04327_ _04329_ u_cpu.cpu.ctrl.o_ibus_adr\[24\]
+ _04337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_83_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05548__A2 _02126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08763_ _04298_ _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05975_ _02486_ _02487_ _02489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07714_ u_cpu.rf_ram.memory\[124\]\[4\] _03553_ _03558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04926_ _01506_ _01510_ _01481_ _01511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08498__A1 _02265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08694_ u_arbiter.i_wb_cpu_dbus_adr\[4\] u_arbiter.i_wb_cpu_dbus_adr\[5\] _04257_
+ _04260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04857_ u_cpu.cpu.decode.opcode\[2\] _01444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07645_ _03506_ _03513_ _03519_ _00706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11114__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07576_ u_cpu.rf_ram.memory\[130\]\[2\] _03475_ _03478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06527_ _02681_ _02872_ _02874_ _00233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09315_ u_cpu.rf_ram.memory\[69\]\[7\] _04613_ _04621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05159__S1 _01509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09246_ _04582_ _04583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06458_ _02687_ _02829_ _02834_ _00204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07473__A2 _03415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05484__A1 _01621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05409_ _01638_ _01989_ _01534_ _01990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09177_ u_cpu.rf_ram.memory\[99\]\[1\] _04543_ _04545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06389_ _02793_ _02794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08128_ _03705_ _03790_ _03797_ _00912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07225__A2 _03277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08422__A1 _02290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08973__A2 _04425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08059_ _02780_ _02965_ _03759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05331__S1 _01509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05787__A2 u_cpu.cpu.ctrl.i_iscomp vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11070_ u_cpu.cpu.o_wdata0 io_in[4] u_cpu.rf_ram_if.wdata0_r\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08710__S _04257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10021_ _00415_ io_in[4] u_cpu.rf_ram.memory\[61\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06736__A1 _02891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05539__A2 _02117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05354__B _01558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09150__A2 _04523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05073__C _01486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10923_ _01292_ io_in[4] u_cpu.rf_ram.memory\[59\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07161__A1 _03110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10854_ _01223_ io_in[4] u_cpu.rf_ram.memory\[79\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05711__A2 _02286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09340__I _02666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10785_ _01154_ io_in[4] u_cpu.rf_ram.memory\[96\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07464__A2 _03415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05475__A1 _01464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10631__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08413__A1 _03914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07216__A2 _03267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05322__S1 _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06975__A1 _03104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10781__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10219_ _00605_ io_in[4] u_cpu.rf_ram.memory\[39\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10011__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11137__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05760_ _02316_ _02335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_36_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09141__A2 _04523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05691_ u_arbiter.i_wb_cpu_dbus_we _02266_ u_cpu.cpu.immdec.imm24_20\[0\] _02268_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_36_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07430_ u_cpu.rf_ram.memory\[137\]\[1\] _03395_ _03397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10161__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07361_ _03312_ _03355_ _03358_ _00583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06312_ _02637_ _02745_ _02747_ _00145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09100_ _04501_ _01180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07455__A2 _03405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07292_ u_cpu.rf_ram.memory\[72\]\[5\] _03308_ _03319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09031_ u_cpu.rf_ram.memory\[96\]\[1\] _04463_ _04465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05010__S0 _01496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06243_ u_cpu.rf_ram.memory\[81\]\[7\] _02697_ _02705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08404__A1 _03901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07207__A2 _03267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06174_ _02606_ u_cpu.rf_ram_if.wdata1_r\[5\] _02654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_116_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05125_ _01597_ _01708_ _01600_ _01709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05313__S1 _01500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05769__A2 _02277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09933_ _00327_ io_in[4] u_cpu.rf_ram.memory\[76\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05056_ _01522_ _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09864_ _00258_ io_in[4] u_cpu.rf_ram_if.rcnt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06718__A1 _02891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__04997__C _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08815_ u_cpu.cpu.ctrl.o_ibus_adr\[15\] _04327_ _04311_ u_cpu.cpu.ctrl.o_ibus_adr\[16\]
+ _04328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09795_ _00189_ io_in[4] u_cpu.rf_ram.memory\[45\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05174__B _01518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08746_ u_arbiter.i_wb_cpu_dbus_adr\[30\] u_arbiter.i_wb_cpu_dbus_adr\[31\] _02335_
+ _04286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05958_ _02456_ _02474_ _02475_ _00062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_39_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09132__A2 _04513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10504__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04909_ u_cpu.raddr\[0\] _01494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_54_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08677_ u_cpu.rf_ram.memory\[31\]\[3\] _04247_ _04251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05889_ _02430_ _00035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_42_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07143__A1 _03110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07628_ _03508_ _03496_ _03509_ _00699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07694__A2 _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07559_ _03312_ _03465_ _03468_ _00671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10654__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10570_ _00943_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07446__A2 _03405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08932__C _03969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09229_ u_cpu.rf_ram.memory\[106\]\[0\] _04573_ _04574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05552__S1 _01594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09199__A2 _04553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05209__A1 _01490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08946__A2 _03910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05304__S1 _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06957__A1 _03104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11122_ _00053_ io_in[0] u_scanchain_local.module_data_in\[34\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11053_ _01422_ io_in[4] u_cpu.rf_ram.memory\[89\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10034__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06709__A1 u_cpu.rf_ram.memory\[139\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10004_ _00398_ io_in[4] u_cpu.rf_ram.memory\[63\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09371__A2 _04651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06185__A2 _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09123__A2 _04513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10184__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10906_ _01275_ io_in[4] u_cpu.rf_ram.memory\[69\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07685__A2 _03533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10837_ _01206_ io_in[4] u_cpu.rf_ram.memory\[104\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05531__C _01560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08634__A1 _04013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07437__A2 _03395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10768_ _01137_ io_in[4] u_cpu.rf_ram.memory\[94\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10699_ _01069_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05543__S1 _01524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06930_ u_cpu.rf_ram.memory\[29\]\[7\] _03100_ _03115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06861_ _02889_ _03069_ _03073_ _00368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10527__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08600_ _04173_ _04052_ _04111_ _04190_ _04191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_95_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05812_ _02272_ u_cpu.rf_ram_if.rdata1\[6\] _02380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09580_ u_cpu.rf_ram.memory\[25\]\[7\] _04772_ _04780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06792_ _02893_ _03028_ _03034_ _00338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09114__A2 _04503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08531_ _04127_ _04129_ _04053_ _04130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05743_ _01444_ _02265_ _02318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07125__A1 _03110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10677__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05674_ u_cpu.rf_ram.memory\[140\]\[7\] u_cpu.rf_ram.memory\[141\]\[7\] u_cpu.rf_ram.memory\[142\]\[7\]
+ u_cpu.rf_ram.memory\[143\]\[7\] _01523_ _01525_ _02252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08462_ _03955_ _04068_ _04070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07676__A2 _03533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07413_ _03310_ _03385_ _03387_ _00606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08393_ _04000_ _03931_ _04013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07344_ u_cpu.rf_ram.memory\[70\]\[3\] _03345_ _03349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08625__A1 _03923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07428__A2 _03395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08525__S _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05013__I _01495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07275_ _02768_ _02954_ _03307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05534__S1 _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09014_ _04438_ _04453_ _04455_ _01140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06226_ _02614_ _02672_ _02695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_128_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08928__A2 _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05169__B _01482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06157_ _02611_ u_cpu.rf_ram_if.wdata0_r\[2\] _02639_ _02640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10057__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09050__A1 _02677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06939__A1 _03104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05884__S _02418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05108_ _01512_ _01691_ _01692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05298__S0 _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06088_ _02397_ _02579_ _02580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07600__A2 _03485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09916_ _00310_ io_in[4] u_cpu.rf_ram.memory\[77\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05039_ _01621_ _01623_ _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09353__A2 _04641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09847_ _00241_ io_in[4] u_cpu.rf_ram.memory\[50\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06167__A2 _02647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08994__I _02646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09778_ _00172_ io_in[4] u_cpu.rf_ram.memory\[42\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09105__A2 _04503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05470__S0 _01576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08729_ _04277_ _01033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07667__A2 _03523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10622_ _00995_ io_in[4] u_cpu.cpu.immdec.imm31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07419__A2 _03385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10553_ _00926_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08092__A2 _03770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05525__S1 _01499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10484_ _00857_ io_in[4] u_cpu.rf_ram.memory\[121\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08919__A2 _04381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05850__A1 u_cpu.cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09592__A2 _04782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11105_ _00034_ io_in[0] u_arbiter.i_wb_cpu_rdt\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09842__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11036_ _01405_ io_in[4] u_cpu.rf_ram.memory\[98\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05461__S0 _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07107__A1 _03110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09992__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05542__B _02120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07658__A2 _03523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04937__I _01495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05669__A1 _02227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06330__A2 _02756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05390_ u_cpu.rf_ram.memory\[80\]\[4\] u_cpu.rf_ram.memory\[81\]\[4\] u_cpu.rf_ram.memory\[82\]\[4\]
+ u_cpu.rf_ram.memory\[83\]\[4\] _01544_ _01545_ _01971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_13_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04892__A2 _01452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08083__A2 _03770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09280__A1 _04450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05516__S1 _01532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06094__A1 _02305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07060_ u_cpu.rf_ram.memory\[57\]\[0\] _03187_ _03188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07830__A2 _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06011_ _02418_ u_scanchain_local.module_data_in\[53\] _02398_ u_arbiter.i_wb_cpu_dbus_adr\[16\]
+ _02517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__09032__A1 _04438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06397__A2 _02794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07962_ _03703_ _03693_ _03704_ _00839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09701_ _02927_ _04847_ _01435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09335__A2 _04624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06913_ _03102_ _03100_ _03103_ _00390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06149__A2 _02632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07893_ u_cpu.rf_ram.memory\[35\]\[1\] _03662_ _03664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11157__D _00091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09632_ u_cpu.rf_ram.memory\[98\]\[6\] _04802_ _04809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06844_ u_cpu.rf_ram.memory\[67\]\[4\] _03059_ _03064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07897__A2 _03662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09563_ _04638_ _04762_ _04770_ _01374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06775_ u_cpu.rf_ram.memory\[76\]\[6\] _03018_ _03025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08514_ _04111_ _04112_ _04114_ _03910_ _03966_ _04115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_05726_ _01460_ _02301_ _02302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09494_ u_cpu.cpu.state.genblk1.misalign_trap_sync_r _04724_ _04726_ _04727_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07649__A2 _03513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05204__S0 _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08445_ _03935_ _03974_ _04054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05657_ _01554_ _02234_ _01607_ _02235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_23_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06321__A2 _02745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08376_ _03997_ _03972_ _03998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05588_ u_cpu.rf_ram.memory\[140\]\[6\] u_cpu.rf_ram.memory\[141\]\[6\] u_cpu.rf_ram.memory\[142\]\[6\]
+ u_cpu.rf_ram.memory\[143\]\[6\] _01641_ _01642_ _02167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_20_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09715__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07327_ _03314_ _03335_ _03339_ _00568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08074__A2 _03760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05507__S1 _01509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07258_ u_cpu.rf_ram.memory\[13\]\[0\] _03297_ _03298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07821__A2 _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06209_ u_cpu.rf_ram.memory\[21\]\[2\] _02679_ _02684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07189_ _02637_ _03257_ _03259_ _00510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09574__A2 _04772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09865__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06388__A2 _02782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07585__A1 _03320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05627__B _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10842__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09326__A2 _04624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05346__C _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07888__A2 _03652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10992__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06312__A2 _02745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10222__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10605_ _00978_ io_in[4] u_cpu.cpu.immdec.imm24_20\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08065__A2 _03760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09262__A1 _04450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06193__B _01494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10536_ _00909_ io_in[4] u_cpu.rf_ram.memory\[33\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10372__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05823__A1 _01467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09014__A1 _04438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10467_ _00840_ io_in[4] u_cpu.rf_ram.memory\[120\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06379__A2 _02784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10398_ _00771_ io_in[4] u_cpu.rf_ram.memory\[36\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11019_ _01388_ io_in[4] u_cpu.rf_ram.memory\[24\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04890_ _01448_ _01443_ _01457_ _01477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__07879__A2 _03652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06000__A1 _02402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08567__C _02318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06560_ _02661_ _02895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_64_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05511_ u_cpu.rf_ram.memory\[16\]\[6\] u_cpu.rf_ram.memory\[17\]\[6\] u_cpu.rf_ram.memory\[18\]\[6\]
+ u_cpu.rf_ram.memory\[19\]\[6\] _01508_ _01509_ _02090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09738__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06491_ u_cpu.rf_ram.memory\[43\]\[2\] _02851_ _02854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06303__A2 _02733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05442_ _01463_ _02021_ _01558_ _02022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08230_ _03872_ _03873_ _00938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10715__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05373_ u_cpu.rf_ram.memory\[104\]\[4\] u_cpu.rf_ram.memory\[105\]\[4\] u_cpu.rf_ram.memory\[106\]\[4\]
+ u_cpu.rf_ram.memory\[107\]\[4\] _01555_ _01531_ _01954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08161_ _02416_ _03822_ _03825_ _00917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08056__A2 _03750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07112_ _02827_ _03037_ _03216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08092_ _03705_ _03770_ _03777_ _00896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09888__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07043_ _03098_ _03177_ _03178_ _00445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09005__A1 _04448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10865__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09556__A2 _04762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07567__A1 _03320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05447__B _01480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08994_ _02646_ _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09308__A2 _04613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07945_ _03692_ _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08516__B1 _04106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06790__A2 _03028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08516__C2 _04009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07876_ _03498_ _03652_ _03654_ _00803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08477__C _03912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09615_ _02691_ _04792_ _04799_ _01397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06827_ _02891_ _03049_ _03054_ _00353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10245__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09546_ _02677_ _02780_ _04761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06758_ _02895_ _03008_ _03015_ _00323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05709_ _01441_ _02285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09477_ u_cpu.rf_ram.memory\[88\]\[3\] _04711_ _04715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09492__A1 u_cpu.cpu.decode.op21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06689_ _02695_ _02976_ _02977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08428_ _03695_ _04041_ _04043_ _00966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10395__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04856__A2 u_cpu.cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08047__A2 _03750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09244__A1 _04450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08359_ _02305_ _03956_ _03940_ _03959_ _03983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_137_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05805__A1 _02273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10321_ _00707_ io_in[4] u_cpu.rf_ram.memory\[128\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10252_ _00638_ io_in[4] u_cpu.rf_ram.memory\[135\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10183_ _00569_ io_in[4] u_cpu.rf_ram.memory\[71\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06230__A1 _02669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11020__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06781__A2 _03028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08522__A3 _04051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06533__A2 _02872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10738__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08286__A2 u_arbiter.i_wb_cpu_rdt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08038__A2 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10888__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07797__A1 u_cpu.cpu.state.o_cnt_r\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10519_ _00892_ io_in[4] u_cpu.rf_ram.memory\[115\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09538__A2 _04752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10118__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07549__A1 _03320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08210__A2 _03835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05991_ _02389_ u_scanchain_local.module_data_in\[48\] _02398_ u_arbiter.i_wb_cpu_dbus_adr\[11\]
+ _02501_ _02502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_66_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06772__A2 _03018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07730_ u_cpu.rf_ram.memory\[123\]\[3\] _03563_ _03567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10268__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04942_ _01493_ _01526_ _01527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07661_ _03504_ _03523_ _03528_ _00713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04873_ u_cpu.cpu.state.genblk1.misalign_trap_sync_r _01459_ _01460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06524__A2 _02872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07721__A1 _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06098__B _02305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09400_ _04622_ _04671_ _04672_ _01309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06612_ _01635_ _02930_ _02933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_81_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07592_ u_cpu.rf_ram.memory\[12\]\[1\] _03485_ _03487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09331_ _02651_ _04632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06543_ u_cpu.rf_ram.memory\[50\]\[0\] _02883_ _02884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09474__A1 _04626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09262_ _04450_ _04583_ _04591_ _01252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06474_ u_cpu.rf_ram.memory\[41\]\[3\] _02840_ _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08213_ u_arbiter.i_wb_cpu_dbus_dat\[19\] _03808_ _03862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05425_ _01998_ _02000_ _02002_ _02004_ _01486_ _02005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_21_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09193_ u_cpu.rf_ram.memory\[79\]\[0\] _04553_ _04554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09226__A1 _04450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08029__A2 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09077__I1 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08144_ u_arbiter.i_wb_cpu_dbus_dat\[0\] u_arbiter.i_wb_cpu_dbus_dat\[1\] _02915_
+ _03811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05356_ u_cpu.rf_ram.memory\[60\]\[4\] u_cpu.rf_ram.memory\[61\]\[4\] u_cpu.rf_ram.memory\[62\]\[4\]
+ u_cpu.rf_ram.memory\[63\]\[4\] _01496_ _01594_ _01937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_107_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05287_ _01862_ _01864_ _01866_ _01868_ _01560_ _01869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_119_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08075_ u_cpu.rf_ram.memory\[122\]\[7\] _03760_ _03768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07026_ u_cpu.rf_ram.memory\[5\]\[1\] _03167_ _03169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06460__A1 _02689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11043__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08201__A2 _03835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05646__S0 _01576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08977_ u_cpu.rf_ram.memory\[97\]\[5\] _04425_ _04431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06763__A2 _03018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09903__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07928_ _03494_ _03682_ _03683_ _00826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07859_ _03639_ _03641_ _03642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_29_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06515__A2 _02861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08760__I0 _02355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10870_ _01239_ io_in[4] u_cpu.rf_ram.memory\[106\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08708__S _04257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09529_ _04751_ _04752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08512__I0 u_arbiter.i_wb_cpu_rdt\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07779__A1 _03494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08440__A2 _04041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10304_ _00690_ io_in[4] u_cpu.rf_ram.memory\[12\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10235_ _00621_ io_in[4] u_cpu.rf_ram.memory\[49\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10410__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05637__S0 _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10166_ _00552_ io_in[4] u_cpu.rf_ram.memory\[72\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06754__A2 _03008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05962__B1 _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10097_ _00491_ io_in[4] u_cpu.rf_ram.memory\[53\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10560__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07703__A1 _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06506__A2 _02861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05190__A1 _01492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09456__A1 _04626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08259__A2 _03885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10999_ _01368_ io_in[4] u_cpu.rf_ram.memory\[26\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05550__B _01480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04945__I _01529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09208__A1 _04450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05868__I1 u_arbiter.i_wb_cpu_dbus_dat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05210_ u_cpu.rf_ram.memory\[92\]\[2\] u_cpu.rf_ram.memory\[93\]\[2\] u_cpu.rf_ram.memory\[94\]\[2\]
+ u_cpu.rf_ram.memory\[95\]\[2\] _01562_ _01563_ _01793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_50_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06190_ u_cpu.rf_ram.memory\[82\]\[7\] _02628_ _02668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11066__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05141_ _01705_ _01724_ _01471_ _01725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08431__A2 _04041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05072_ _01506_ _01655_ _01519_ _01656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_131_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06993__A2 _03147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08900_ u_cpu.rf_ram.memory\[2\]\[4\] _04371_ _04376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09926__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09880_ _00274_ io_in[4] u_cpu.rf_ram.memory\[17\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10090__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08831_ _04336_ _01076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07942__A1 _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10903__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06745__A2 _03008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08762_ _02677_ _02766_ _04298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05953__B1 _02398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05974_ _02486_ _02487_ _02488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07713_ _03502_ _03553_ _03557_ _00736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_04925_ u_cpu.rf_ram.memory\[24\]\[0\] u_cpu.rf_ram.memory\[25\]\[0\] u_cpu.rf_ram.memory\[26\]\[0\]
+ u_cpu.rf_ram.memory\[27\]\[0\] _01508_ _01509_ _01510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08693_ _04259_ _01015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09695__A1 _02273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07644_ u_cpu.rf_ram.memory\[128\]\[5\] _03513_ _03519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04856_ _01441_ u_cpu.cpu.bne_or_bge _01442_ _01443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__07170__A2 _03247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07575_ _03310_ _03475_ _03477_ _00678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05181__A1 _01464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09314_ _04448_ _04613_ _04620_ _01275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06526_ u_cpu.rf_ram.memory\[47\]\[1\] _02872_ _02874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09245_ _02849_ _04349_ _04582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06457_ u_cpu.rf_ram.memory\[51\]\[4\] _02829_ _02834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06681__A1 _02891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05484__A2 _02063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05408_ u_cpu.rf_ram.memory\[140\]\[4\] u_cpu.rf_ram.memory\[141\]\[4\] u_cpu.rf_ram.memory\[142\]\[4\]
+ u_cpu.rf_ram.memory\[143\]\[4\] _01634_ _01635_ _01989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_119_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09176_ _04434_ _04543_ _04544_ _01213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06388_ _02766_ _02782_ _02793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08127_ u_cpu.rf_ram.memory\[33\]\[6\] _03790_ _03797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05339_ _01493_ _01919_ _01920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08422__A2 _03956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10433__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06433__A1 _02683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08058_ _03707_ _03750_ _03758_ _00881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05619__C _01560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06984__A2 _03137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07009_ _03102_ _03157_ _03159_ _00430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08997__I _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04995__A1 _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08186__A1 u_arbiter.i_wb_cpu_dbus_dat\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10020_ _00414_ io_in[4] u_cpu.rf_ram.memory\[61\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10583__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06736__A2 _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11075__D u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10922_ _01291_ io_in[4] u_cpu.rf_ram.memory\[59\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07161__A2 _03237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09438__A1 _04626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10853_ _01222_ io_in[4] u_cpu.rf_ram.memory\[79\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05172__A1 _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05370__B _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10784_ _01153_ io_in[4] u_cpu.rf_ram.memory\[96\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08110__A1 _03705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11089__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08661__A2 _04237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05475__A2 _02054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09949__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08413__A2 _03938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09068__I _02910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06424__A1 _02693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10926__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06975__A2 _03137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10218_ _00604_ io_in[4] u_cpu.rf_ram.memory\[138\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06727__A2 _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07924__A1 _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10149_ _00535_ io_in[4] u_cpu.rf_ram.memory\[140\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06220__I _02661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09677__A1 _04626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05690_ u_arbiter.i_wb_cpu_dbus_we _02264_ _02266_ _02267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_35_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07152__A2 _03237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10306__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05163__A1 _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07360_ u_cpu.rf_ram.memory\[143\]\[2\] _03355_ _03358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06311_ u_cpu.rf_ram.memory\[7\]\[1\] _02745_ _02747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07291_ _02656_ _03318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10456__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09030_ _04434_ _04463_ _04464_ _01147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05010__S1 _01594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06242_ _02691_ _02697_ _02704_ _00118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06173_ _02628_ _02652_ _02653_ _00100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05218__A2 _01796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05124_ u_cpu.rf_ram.memory\[88\]\[1\] u_cpu.rf_ram.memory\[89\]\[1\] u_cpu.rf_ram.memory\[90\]\[1\]
+ u_cpu.rf_ram.memory\[91\]\[1\] _01598_ _01556_ _01708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__05069__I2 u_cpu.rf_ram.memory\[22\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06966__A2 _03127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09932_ _00326_ io_in[4] u_cpu.rf_ram.memory\[76\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05055_ _01638_ _01639_ _01534_ _01640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09863_ _00257_ io_in[4] u_cpu.rf_ram_if.rcnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06718__A2 _02988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08814_ _04308_ _04327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09794_ _00188_ io_in[4] u_cpu.rf_ram.memory\[45\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08745_ _04285_ _01041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_73_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05957_ _02389_ u_scanchain_local.module_data_in\[41\] _02398_ u_arbiter.i_wb_cpu_dbus_adr\[4\]
+ _02475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04908_ _01464_ _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08676_ _03697_ _04247_ _04250_ _01007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05888_ u_arbiter.i_wb_cpu_rdt\[15\] u_arbiter.i_wb_cpu_dbus_dat\[12\] _02418_ _02430_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08340__A1 _02911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07143__A2 _03227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08485__C _04031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07627_ u_cpu.rf_ram.memory\[22\]\[6\] _03496_ _03509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05154__A1 _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05190__B _01772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04901__A1 u_cpu.cpu.immdec.imm24_20\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07558_ u_cpu.rf_ram.memory\[131\]\[2\] _03465_ _03468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06509_ u_cpu.rf_ram.memory\[48\]\[2\] _02861_ _02864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07489_ _03314_ _03425_ _03429_ _00640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09089__S _04485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09228_ _04572_ _04573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06654__A1 _02881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10949__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09159_ u_cpu.rf_ram.memory\[104\]\[1\] _04533_ _04535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05209__A2 _01782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06957__A2 _03127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11121_ _00052_ io_in[0] u_arbiter.i_wb_cpu_rdt\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04968__A1 _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08159__A1 _02915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11052_ _01421_ io_in[4] u_cpu.rf_ram.memory\[89\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06709__A2 _02988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07906__A1 _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10003_ _00397_ io_in[4] u_cpu.rf_ram.memory\[63\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07382__A2 _03365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10329__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05393__A1 _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09659__A1 _04626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08331__A1 _02466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07134__A2 _03227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10905_ _01274_ io_in[4] u_cpu.rf_ram.memory\[69\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05145__A1 _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08882__A2 _04361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10479__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10836_ _01205_ io_in[4] u_cpu.rf_ram.memory\[104\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06893__A1 _02885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10767_ _01136_ io_in[4] u_cpu.rf_ram.memory\[94\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09771__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06645__A1 _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10698_ _01068_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05999__A3 _02499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06948__A2 _03117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11104__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05275__B _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06860_ u_cpu.rf_ram.memory\[66\]\[3\] _03069_ _03073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05811_ _02273_ u_cpu.rf_ram.rdata\[6\] _02379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06791_ u_cpu.rf_ram.memory\[75\]\[5\] _03028_ _03034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08530_ _04055_ _04128_ _04129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05742_ _02306_ _02316_ _02317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_36_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07125__A2 _03217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08461_ _03896_ _04068_ _04069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__05136__A1 _01621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05673_ _01638_ _02250_ _01482_ _02251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_63_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07412_ u_cpu.rf_ram.memory\[39\]\[1\] _03385_ _03387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08392_ _03899_ _03917_ _03962_ _04012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_50_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07343_ _03312_ _03345_ _03348_ _00575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08625__A2 _04052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07274_ _02631_ _03306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09013_ u_cpu.rf_ram.memory\[95\]\[1\] _04453_ _04455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06225_ _02693_ _02679_ _02694_ _00111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08389__A1 _03895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06156_ _02606_ u_cpu.rf_ram_if.wdata1_r\[2\] _02639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09050__A2 _02814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06939__A2 _03117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05107_ u_cpu.rf_ram.memory\[108\]\[1\] u_cpu.rf_ram.memory\[109\]\[1\] u_cpu.rf_ram.memory\[110\]\[1\]
+ u_cpu.rf_ram.memory\[111\]\[1\] _01551_ _01524_ _01691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_132_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07061__A1 _03098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05298__S1 _01563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06087_ u_cpu.cpu.ctrl.o_ibus_adr\[30\] _02577_ _02579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09915_ _00309_ io_in[4] u_cpu.rf_ram.memory\[77\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05038_ u_cpu.rf_ram.memory\[64\]\[0\] u_cpu.rf_ram.memory\[65\]\[0\] u_cpu.rf_ram.memory\[66\]\[0\]
+ u_cpu.rf_ram.memory\[67\]\[0\] _01522_ _01622_ _01623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_99_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09846_ _00240_ io_in[4] u_cpu.rf_ram.memory\[50\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07364__A2 _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09777_ _00171_ io_in[4] u_cpu.rf_ram.memory\[42\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06989_ _03098_ _03147_ _03148_ _00421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08728_ u_arbiter.i_wb_cpu_dbus_adr\[21\] u_arbiter.i_wb_cpu_dbus_adr\[22\] _02335_
+ _04277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05470__S1 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10621__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07116__A2 _03217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05127__A1 _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08659_ u_cpu.rf_ram.memory\[32\]\[3\] _04237_ _04241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09794__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08864__A2 _04351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06875__A1 _02885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08716__S _04257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05922__I0 u_arbiter.i_wb_cpu_rdt\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10621_ _00994_ io_in[4] u_cpu.cpu.immdec.imm19_12_20\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10771__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06627__A1 _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10552_ _00925_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10483_ _00856_ io_in[4] u_cpu.rf_ram.memory\[121\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11127__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10001__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05850__A2 _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09041__A2 _04463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11104_ _00033_ io_in[0] u_arbiter.i_wb_cpu_rdt\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10151__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11035_ _01404_ io_in[4] u_cpu.rf_ram.memory\[98\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05095__B _01480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08552__A1 _03969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05366__A1 _01492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05461__S1 _01531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07107__A2 _03207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05913__I0 u_arbiter.i_wb_cpu_rdt\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10819_ _01188_ io_in[4] u_cpu.rf_ram.memory\[101\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04972__S0 _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08607__A2 _03955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09280__A2 _04593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06010_ u_cpu.cpu.ctrl.o_ibus_adr\[16\] _02515_ _02516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_12_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09032__A2 _04463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07043__A1 _03098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08240__B1 _03829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07594__A2 _03485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07961_ u_cpu.rf_ram.memory\[120\]\[5\] _03693_ _03704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09700_ _02912_ _04846_ _04847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06912_ u_cpu.rf_ram.memory\[29\]\[1\] _03100_ _03103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07892_ _03494_ _03662_ _03663_ _00810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10644__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08543__A1 _04009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07346__A2 _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09631_ _04634_ _04802_ _04808_ _01404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08543__B2 _03955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06843_ _02889_ _03059_ _03063_ _00360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05357__A1 _01464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09562_ u_cpu.rf_ram.memory\[26\]\[7\] _04762_ _04770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06774_ _02893_ _03018_ _03024_ _00330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08513_ _03932_ _04051_ _04113_ _03909_ _04114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05725_ _02282_ _02284_ _02287_ _02288_ _02300_ _02301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_70_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10794__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09493_ u_cpu.cpu.genblk3.csr.o_new_irq _04725_ _04726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05452__C _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08846__A2 _04327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05204__S1 _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06857__A1 _02885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08444_ _04000_ _04052_ _03915_ _04053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05656_ u_cpu.rf_ram.memory\[84\]\[7\] u_cpu.rf_ram.memory\[85\]\[7\] u_cpu.rf_ram.memory\[86\]\[7\]
+ u_cpu.rf_ram.memory\[87\]\[7\] _01507_ _01605_ _02234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_23_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08375_ _03974_ _03947_ _03997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05587_ _01493_ _02165_ _02166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10024__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06609__A1 _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07326_ u_cpu.rf_ram.memory\[71\]\[3\] _03335_ _03339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09271__A2 _04593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07257_ _03296_ _03297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05895__S _02431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06208_ _02641_ _02683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05832__A2 u_cpu.cpu.state.o_cnt_r\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09023__A2 _04453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07188_ u_cpu.rf_ram.memory\[15\]\[1\] _03257_ _03259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10174__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06139_ _02608_ _02623_ _02624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08782__A1 _02395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07585__A2 _03475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05596__A1 _01506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08534__A1 _03906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09829_ _00223_ io_in[4] u_cpu.rf_ram.memory\[43\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05348__A1 _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05643__B _01558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11083__D u_cpu.rf_ram_if.wdata1_r\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08954__B _04031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10604_ _00977_ io_in[4] u_cpu.cpu.immdec.imm24_20\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09262__A2 _04583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10517__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06076__A2 _02562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07273__A1 _02667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10535_ _00908_ io_in[4] u_cpu.rf_ram.memory\[33\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10466_ _00839_ io_in[4] u_cpu.rf_ram.memory\[120\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09014__A2 _04453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07025__A1 _02632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10397_ _00770_ io_in[4] u_cpu.rf_ram.memory\[36\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10667__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08773__A1 _03701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07576__A2 _03475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05131__S0 _01522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05587__A1 _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07328__A2 _03335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11018_ _01387_ io_in[4] u_cpu.rf_ram.memory\[24\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05339__A1 _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08828__A2 _04327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10047__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05510_ _01513_ _02088_ _02089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06839__A1 _02885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06490_ _02681_ _02851_ _02853_ _00217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07500__A2 _03435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05441_ u_cpu.rf_ram.memory\[44\]\[5\] u_cpu.rf_ram.memory\[45\]\[5\] u_cpu.rf_ram.memory\[46\]\[5\]
+ u_cpu.rf_ram.memory\[47\]\[5\] _01555_ _01531_ _02021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_53_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05362__I1 u_cpu.rf_ram.memory\[49\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08160_ u_arbiter.i_wb_cpu_dbus_dat\[3\] _03818_ _03824_ _03802_ _03807_ _03825_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_05372_ _01512_ _01952_ _01953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09253__A2 _04583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10197__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07111_ _03114_ _03207_ _03215_ _00476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08091_ u_cpu.rf_ram.memory\[115\]\[6\] _03770_ _03777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05814__A2 _01467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07042_ u_cpu.rf_ram.memory\[58\]\[0\] _03177_ _03178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09005__A2 _04436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07567__A2 _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08993_ _04440_ _04436_ _04441_ _01133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05122__S0 _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05578__A1 _01617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07944_ _02954_ _02965_ _03692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07875_ u_cpu.rf_ram.memory\[92\]\[1\] _03652_ _03654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09614_ u_cpu.rf_ram.memory\[0\]\[6\] _04792_ _04799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06826_ u_cpu.rf_ram.memory\[68\]\[4\] _03049_ _03054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09545_ _04638_ _04752_ _04760_ _01366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06757_ u_cpu.rf_ram.memory\[74\]\[6\] _03008_ _03015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05708_ _01442_ u_cpu.cpu.alu.i_rs1 _02283_ _02284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09476_ _04628_ _04711_ _04714_ _01343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06688_ _02608_ _02622_ _02976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09492__A2 _01443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08427_ u_cpu.rf_ram.memory\[114\]\[1\] _04041_ _04043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05639_ _02210_ _02212_ _02214_ _02216_ _01560_ _02217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08358_ _02400_ _03956_ _03982_ _00957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__04856__A3 _01442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09832__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09244__A2 _04573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07255__A1 _03114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07309_ _03314_ _03325_ _03329_ _00560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08289_ _02909_ u_arbiter.i_wb_cpu_rdt\[13\] _03916_ _03917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09097__S _04485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10320_ _00706_ io_in[4] u_cpu.rf_ram.memory\[128\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07007__A1 _03098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09982__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10251_ _00637_ io_in[4] u_cpu.rf_ram.memory\[135\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05638__B _01480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08755__A1 _02596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07558__A2 _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05569__A1 _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10182_ _00568_ io_in[4] u_cpu.rf_ram.memory\[71\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06230__A2 _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08507__A1 _03944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09180__A1 _04440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07730__A2 _03563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09483__A2 _04711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06297__A2 _02733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09235__A2 _04573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10518_ _00891_ io_in[4] u_cpu.rf_ram.memory\[115\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10449_ _00822_ io_in[4] u_cpu.rf_ram.memory\[34\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07549__A2 _03455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06223__I _02666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05267__C _01560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06221__A2 _02679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05990_ _02499_ _02500_ _02456_ _02501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04941_ u_cpu.rf_ram.memory\[4\]\[0\] u_cpu.rf_ram.memory\[5\]\[0\] u_cpu.rf_ram.memory\[6\]\[0\]
+ u_cpu.rf_ram.memory\[7\]\[0\] _01523_ _01525_ _01526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_66_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09705__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07660_ u_cpu.rf_ram.memory\[127\]\[4\] _03523_ _03528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04872_ u_cpu.cpu.decode.op21 _01443_ _01457_ _01458_ _01459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07721__A2 _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06611_ _02932_ _00259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_65_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05732__A1 u_cpu.cpu.genblk3.csr.o_new_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07591_ _02632_ _03485_ _03486_ _00685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_53_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09330_ _04630_ _04624_ _04631_ _01280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06542_ _02882_ _02883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09855__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09474__A2 _04711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09261_ u_cpu.rf_ram.memory\[107\]\[7\] _04583_ _04591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07485__A1 _03310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06473_ _02683_ _02840_ _02843_ _00210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08212_ _03860_ _03861_ _00932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05424_ _01506_ _02003_ _01519_ _02004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_18_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10832__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09192_ _04552_ _04553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09226__A2 _04563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08143_ u_arbiter.i_wb_cpu_dbus_dat\[2\] _02915_ _03810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07237__A1 _03114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05355_ _01929_ _01931_ _01933_ _01935_ _01560_ _01936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_88_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07788__A2 _03593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08074_ _03705_ _03760_ _03767_ _00888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05286_ _01566_ _01867_ _01558_ _01868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05799__A1 _02273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07025_ _02632_ _03167_ _03168_ _00437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10982__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05458__B _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06460__A2 _02829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06212__A2 _02679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05646__S1 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10212__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08976_ _03701_ _04425_ _04430_ _01127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07927_ u_cpu.rf_ram.memory\[117\]\[0\] _03682_ _03683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05971__A1 _02456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09162__A1 _04440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07858_ _02280_ _03640_ _03641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_60_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07712__A2 _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06809_ _02652_ _03039_ _03044_ _00345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10362__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07789_ _03506_ _03593_ _03599_ _00770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_43_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09528_ _02677_ _02849_ _04751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09465__A2 _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08512__I1 u_arbiter.i_wb_cpu_rdt\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09459_ u_cpu.rf_ram.memory\[87\]\[3\] _04701_ _04705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06279__A2 _02719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08724__S _02335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09217__A2 _04563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05582__S0 _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08976__A1 _03701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07779__A2 _03593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10303_ _00689_ io_in[4] u_cpu.rf_ram.memory\[12\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06451__A2 _02829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10234_ _00620_ io_in[4] u_cpu.rf_ram.memory\[137\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09728__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06203__A2 _02679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05637__S1 _01531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10165_ _00551_ io_in[4] u_cpu.rf_ram.memory\[72\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05962__A1 _02403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10096_ _00490_ io_in[4] u_cpu.rf_ram.memory\[53\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10705__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05962__B2 u_arbiter.i_wb_cpu_dbus_adr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09878__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07703__A2 _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10855__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09456__A2 _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10998_ _01367_ io_in[4] u_cpu.rf_ram.memory\[26\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05190__A2 _01744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07467__A1 _03310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09208__A2 _04553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05573__S0 _01507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07219__A1 _03114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05140_ _01492_ _01714_ _01723_ _01724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_7_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06442__A2 _02816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05071_ u_cpu.rf_ram.memory\[16\]\[1\] u_cpu.rf_ram.memory\[17\]\[1\] u_cpu.rf_ram.memory\[18\]\[1\]
+ u_cpu.rf_ram.memory\[19\]\[1\] _01508_ _01509_ _01655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__05278__B _01859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10235__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08589__B _03925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09392__A1 _04634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08195__A2 _03835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08830_ u_cpu.cpu.ctrl.o_ibus_adr\[22\] _04327_ _04329_ u_cpu.cpu.ctrl.o_ibus_adr\[23\]
+ _04336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07942__A2 _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08761_ _04297_ _01045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10385__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05973_ u_cpu.cpu.ctrl.o_ibus_adr\[7\] u_cpu.cpu.ctrl.o_ibus_adr\[6\] u_cpu.cpu.ctrl.o_ibus_adr\[5\]
+ _02476_ _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05953__A1 _02389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09144__A1 _04440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07712_ u_cpu.rf_ram.memory\[124\]\[3\] _03553_ _03557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04924_ _01499_ _01509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08692_ u_arbiter.i_wb_cpu_dbus_adr\[3\] u_arbiter.i_wb_cpu_dbus_adr\[4\] _04257_
+ _04259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_54_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07643_ _03504_ _03513_ _03518_ _00705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05705__A1 _02259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04855_ u_cpu.cpu.csr_d_sel _01442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07574_ u_cpu.rf_ram.memory\[130\]\[1\] _03475_ _03477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09447__A2 _04691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09313_ u_cpu.rf_ram.memory\[69\]\[6\] _04613_ _04620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06525_ _02669_ _02872_ _02873_ _00232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07458__A1 u_cpu.rf_ram.memory\[49\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09244_ _04450_ _04573_ _04581_ _01244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06456_ _02685_ _02829_ _02833_ _00203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05564__S0 _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05032__I _01463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11010__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05407_ _01465_ _01987_ _01988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09175_ u_cpu.rf_ram.memory\[99\]\[0\] _04543_ _04544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06681__A2 _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06387_ _02693_ _02784_ _02792_ _00175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08126_ _03703_ _03790_ _03796_ _00911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05338_ u_cpu.rf_ram.memory\[4\]\[4\] u_cpu.rf_ram.memory\[5\]\[4\] u_cpu.rf_ram.memory\[6\]\[4\]
+ u_cpu.rf_ram.memory\[7\]\[4\] _01523_ _01525_ _01919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__04871__I u_cpu.cpu.genblk3.csr.o_new_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08057_ u_cpu.rf_ram.memory\[112\]\[7\] _03750_ _03758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07630__A1 u_cpu.rf_ram.memory\[22\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06433__A2 _02816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05269_ _01464_ _01850_ _01851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07008_ u_cpu.rf_ram.memory\[19\]\[1\] _03157_ _03159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04995__A2 _01578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10728__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08186__A2 _03835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07933__A2 _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08959_ _03901_ _03919_ _04419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10878__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09686__A2 _04832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07697__A1 _03504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10921_ _01290_ io_in[4] u_cpu.rf_ram.memory\[59\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10852_ _01221_ io_in[4] u_cpu.rf_ram.memory\[79\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09438__A2 _04691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10108__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07449__A1 _03310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10783_ _01152_ io_in[4] u_cpu.rf_ram.memory\[96\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08110__A2 _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06672__A2 _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10258__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08949__A1 _02728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05307__S0 _01522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09610__A2 _04792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07621__A1 u_cpu.rf_ram.memory\[22\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06424__A2 _02805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08177__A2 _03835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09374__A1 _02657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10217_ _00603_ io_in[4] u_cpu.rf_ram.memory\[138\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07924__A2 _03672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10148_ _00534_ io_in[4] u_cpu.rf_ram.memory\[140\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05935__A1 u_arbiter.i_wb_cpu_ibus_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09126__A1 _04440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10079_ _00473_ io_in[4] u_cpu.rf_ram.memory\[55\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09677__A2 _04832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05538__I1 u_cpu.rf_ram.memory\[49\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04956__I _01540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09429__A2 _04681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05163__A2 _01745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11033__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08101__A2 _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06310_ _02632_ _02745_ _02746_ _00144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_31_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07290_ _03316_ _03308_ _03317_ _00553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08591__C _03955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06241_ u_cpu.rf_ram.memory\[81\]\[6\] _02697_ _02704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07860__A1 _02285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06663__A2 _02956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06172_ u_cpu.rf_ram.memory\[82\]\[4\] _02628_ _02653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05123_ _01464_ _01706_ _01707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07612__A1 u_cpu.rf_ram.memory\[22\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06415__A2 _02805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09931_ _00325_ io_in[4] u_cpu.rf_ram.memory\[76\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05054_ u_cpu.rf_ram.memory\[140\]\[0\] u_cpu.rf_ram.memory\[141\]\[0\] u_cpu.rf_ram.memory\[142\]\[0\]
+ u_cpu.rf_ram.memory\[143\]\[0\] _01634_ _01635_ _01639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_98_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05736__B _01444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08412__I0 u_arbiter.i_wb_cpu_rdt\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09862_ _00256_ io_in[4] u_cpu.rf_ram_if.rreq_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06179__A1 _02628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07915__A2 _03672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08813_ _04326_ _01068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09793_ _00187_ io_in[4] u_cpu.rf_ram.memory\[45\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05956_ u_cpu.cpu.ctrl.o_ibus_adr\[4\] _02473_ _02474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08744_ u_arbiter.i_wb_cpu_dbus_adr\[29\] u_arbiter.i_wb_cpu_dbus_adr\[30\] _02335_
+ _04285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_100_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09668__A2 _04822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04907_ _01487_ _01488_ _01492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07679__A1 _03504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08675_ u_cpu.rf_ram.memory\[31\]\[2\] _04247_ _04250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05887_ _02429_ _00034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_54_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05471__B _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08340__A2 _03965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07626_ _02661_ _03508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06351__A1 _02669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07557_ _03310_ _03465_ _03467_ _00670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10400__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06508_ _02681_ _02861_ _02863_ _00225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07488_ u_cpu.rf_ram.memory\[135\]\[3\] _03425_ _03429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09227_ _02780_ _04349_ _04572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06654__A2 _02956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06439_ _02689_ _02816_ _02822_ _00197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07851__A1 _01444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09158_ _04434_ _04533_ _04534_ _01205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08109_ u_cpu.rf_ram.memory\[116\]\[6\] _03780_ _03787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10550__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05209__A3 _01791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07603__A1 _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08800__B1 _04311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09089_ u_arbiter.i_wb_cpu_rdt\[26\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[10\]
+ _04485_ _04496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_107_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11120_ _00051_ io_in[0] u_arbiter.i_wb_cpu_rdt\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05090__A1 _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09356__A1 _04634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11051_ _01420_ io_in[4] u_cpu.rf_ram.memory\[89\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07906__A2 _03662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10002_ _00396_ io_in[4] u_cpu.rf_ram.memory\[29\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09108__A1 _04440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05393__A2 _01973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09659__A2 _04822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11056__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08331__A2 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10904_ _01273_ io_in[4] u_cpu.rf_ram.memory\[69\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05145__A2 _01728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10835_ _01204_ io_in[4] u_cpu.rf_ram.memory\[103\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06893__A2 _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09916__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10080__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08095__A1 _02717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10766_ _01135_ io_in[4] u_cpu.rf_ram.memory\[94\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07842__A1 _03502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06645__A2 _02945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10697_ _01067_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09595__A1 _04634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07070__A2 _03187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05081__A1 _01513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05810_ _02272_ _02377_ _02378_ _00019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_67_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08570__A2 _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06790_ _02891_ _03028_ _03033_ _00337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06581__A1 _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05741_ _02308_ _02312_ _02315_ u_cpu.cpu.state.stage_two_req _02316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_94_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05291__B _01600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10423__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08460_ _02265_ _02400_ _01446_ _02259_ _04068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_05672_ u_cpu.rf_ram.memory\[132\]\[7\] u_cpu.rf_ram.memory\[133\]\[7\] u_cpu.rf_ram.memory\[134\]\[7\]
+ u_cpu.rf_ram.memory\[135\]\[7\] _01634_ _01635_ _02250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06333__A1 _02683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07411_ _03306_ _03385_ _03386_ _00605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08391_ _03936_ _03949_ _03919_ _03899_ _03938_ _04011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__06884__A2 _03079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07342_ u_cpu.rf_ram.memory\[70\]\[2\] _03345_ _03348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08086__A1 _03699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10573__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07833__A1 _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06636__A2 _02945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07273_ _02667_ _03297_ _03305_ _00548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_136_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09012_ _04434_ _04453_ _04454_ _01139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06224_ u_cpu.rf_ram.memory\[21\]\[7\] _02679_ _02694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08389__A2 _03965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06155_ _02628_ _02637_ _02638_ _00097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05106_ _01548_ _01689_ _01579_ _01690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_117_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06086_ u_cpu.cpu.ctrl.o_ibus_adr\[30\] _02577_ _02578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07061__A2 _03187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05072__A1 _01506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09914_ _00308_ io_in[4] u_cpu.rf_ram.memory\[139\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05037_ _01499_ _01622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08010__A1 _02637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09845_ _00239_ io_in[4] u_cpu.rf_ram.memory\[47\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11079__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09776_ _00170_ io_in[4] u_cpu.rf_ram.memory\[42\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05375__A2 _01951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06988_ u_cpu.rf_ram.memory\[60\]\[0\] _03147_ _03148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08727_ _04276_ _01032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_73_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05939_ _02458_ _02459_ _00058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09939__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05127__A2 _01710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06324__A1 _02667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08658_ _03697_ _04237_ _04240_ _00999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07609_ u_cpu.rf_ram.memory\[22\]\[0\] _03496_ _03497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06875__A2 _03079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10916__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05922__I1 u_arbiter.i_wb_cpu_dbus_dat\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08589_ _04178_ _04180_ _03925_ _04181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08077__A1 _02825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10620_ _00993_ io_in[4] u_cpu.cpu.immdec.imm19_12_20\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07824__A1 _03502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06627__A2 _02935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10551_ _00924_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10482_ _00855_ io_in[4] u_cpu.rf_ram.memory\[121\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08732__S _02335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09577__A1 _04634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07052__A2 _03177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11103_ _00032_ io_in[0] u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05063__A1 _01633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11034_ _01403_ io_in[4] u_cpu.rf_ram.memory\[98\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10446__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05890__I _02388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05366__A2 _01918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10596__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06866__A2 _03069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05913__I1 u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08068__A1 _03699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10818_ _01187_ io_in[4] u_cpu.rf_ram.memory\[101\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__04972__S1 _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06079__B1 _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07815__A1 _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06618__A2 _02935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10749_ _01118_ io_in[4] u_cpu.cpu.immdec.imm11_7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08240__A1 u_arbiter.i_wb_cpu_rdt\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07043__A2 _03177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05286__B _01558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07960_ _02656_ _03703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06911_ _02636_ _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07891_ u_cpu.rf_ram.memory\[35\]\[0\] _03662_ _03663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06003__B1 _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09630_ u_cpu.rf_ram.memory\[98\]\[5\] _04802_ _04808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06842_ u_cpu.rf_ram.memory\[67\]\[3\] _03059_ _03063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05357__A2 _01937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09561_ _04636_ _04762_ _04769_ _01373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06773_ u_cpu.rf_ram.memory\[76\]\[5\] _03018_ _03024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10939__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08512_ u_arbiter.i_wb_cpu_rdt\[27\] u_arbiter.i_wb_cpu_rdt\[11\] _02466_ _04113_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05724_ _02289_ _02276_ _02294_ u_cpu.cpu.genblk3.csr.mstatus_mie _02299_ _02300_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_64_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09492_ u_cpu.cpu.decode.op21 _01443_ _01457_ _04725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_82_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05655_ _01602_ _02232_ _02233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06857__A2 _03069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08443_ _03917_ _04051_ _04052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04868__A1 u_cpu.cpu.decode.op21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08059__A1 _02780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08374_ _02909_ u_arbiter.i_wb_cpu_rdt\[10\] _03995_ _03996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05586_ u_cpu.rf_ram.memory\[136\]\[6\] u_cpu.rf_ram.memory\[137\]\[6\] u_cpu.rf_ram.memory\[138\]\[6\]
+ u_cpu.rf_ram.memory\[139\]\[6\] _01523_ _01642_ _02165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_20_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07325_ _03312_ _03335_ _03338_ _00567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06609__A2 _02929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06136__I u_cpu.cpu.immdec.imm11_7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07256_ _02731_ _02803_ _03296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10319__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09559__A1 _04634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05293__A1 _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06207_ _02681_ _02679_ _02682_ _00105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07187_ _02632_ _03257_ _03258_ _00509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05832__A3 u_cpu.cpu.state.o_cnt_r\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06138_ _02621_ _02622_ _02623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08231__A1 _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07034__A2 _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05045__A1 _01512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08782__A2 _02599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06069_ _02402_ u_scanchain_local.module_data_in\[63\] _02478_ u_arbiter.i_wb_cpu_dbus_adr\[26\]
+ _02565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_132_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10469__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05596__A2 _02173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09761__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09828_ _00222_ io_in[4] u_cpu.rf_ram.memory\[43\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09759_ _00153_ io_in[4] u_cpu.rf_ram.memory\[80\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08298__A1 _03922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06848__A2 _03059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04859__A1 _01444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10603_ _00976_ io_in[4] u_cpu.cpu.immdec.imm24_20\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07273__A2 _03297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10534_ _00907_ io_in[4] u_cpu.rf_ram.memory\[33\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05284__A1 _01512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10465_ _00838_ io_in[4] u_cpu.rf_ram.memory\[120\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07025__A2 _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10396_ _00769_ io_in[4] u_cpu.rf_ram.memory\[36\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08773__A2 _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05131__S1 _01622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06784__A1 _02885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11017_ _01386_ io_in[4] u_cpu.rf_ram.memory\[24\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05339__A2 _01919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08289__A1 _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06839__A2 _03059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05440_ _01505_ _02019_ _02020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09089__I0 u_arbiter.i_wb_cpu_rdt\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05371_ u_cpu.rf_ram.memory\[108\]\[4\] u_cpu.rf_ram.memory\[109\]\[4\] u_cpu.rf_ram.memory\[110\]\[4\]
+ u_cpu.rf_ram.memory\[111\]\[4\] _01529_ _01500_ _01952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_119_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07110_ u_cpu.rf_ram.memory\[55\]\[7\] _03207_ _03215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08090_ _03703_ _03770_ _03776_ _00895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07264__A2 _03297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08461__A1 _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05275__A1 _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07041_ _03176_ _03177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05795__I _02368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10611__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07016__A2 _03157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08213__A1 u_arbiter.i_wb_cpu_dbus_dat\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05027__A1 _01464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09784__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08764__A2 _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08992_ u_cpu.rf_ram.memory\[94\]\[2\] _04436_ _04441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05122__S1 _01563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07943_ _02631_ _03691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10761__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07874_ _03494_ _03652_ _03653_ _00802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06527__A1 _02681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09613_ _02689_ _04792_ _04798_ _01396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_95_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06825_ _02889_ _03049_ _03053_ _00352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05463__C _01560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09544_ u_cpu.rf_ram.memory\[27\]\[7\] _04752_ _04760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11117__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06756_ _02893_ _03008_ _03014_ _00322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_70_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05707_ _01442_ _01439_ _02283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09475_ u_cpu.rf_ram.memory\[88\]\[2\] _04711_ _04714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06687_ _02897_ _02967_ _02975_ _00292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08426_ _03691_ _04041_ _04042_ _00965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05638_ _01566_ _02215_ _01480_ _02216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_24_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10141__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05569_ _01554_ _02147_ _01607_ _02148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08357_ _03969_ _03978_ _03981_ _03982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07308_ u_cpu.rf_ram.memory\[73\]\[3\] _03325_ _03329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07255__A2 _03287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08288_ _02465_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[13\] _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_137_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05266__A1 _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07239_ _03286_ _03287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10291__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10250_ _00636_ io_in[4] u_cpu.rf_ram.memory\[136\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08204__A1 u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07007__A2 _03157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08755__A2 _02914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10181_ _00567_ io_in[4] u_cpu.rf_ram.memory\[71\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05569__A2 _02147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06766__A1 _02885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08507__A2 _03975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06518__A1 _02691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09180__A2 _04543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07191__A1 _02642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07494__A2 _03425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10634__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08443__A1 _03917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07246__A2 _03287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05257__A1 _01513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10517_ _00890_ io_in[4] u_cpu.rf_ram.memory\[115\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10448_ _00821_ io_in[4] u_cpu.rf_ram.memory\[34\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10784__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10379_ _00752_ io_in[4] u_cpu.rf_ram.memory\[38\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04940_ _01524_ _01525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10014__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04959__I _01495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09171__A2 _04533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04871_ u_cpu.cpu.genblk3.csr.o_new_irq _01458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_66_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06610_ _02912_ _02927_ _02930_ _02931_ _02932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_19_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07590_ u_cpu.rf_ram.memory\[12\]\[0\] _03485_ _03486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_92_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05732__A2 u_cpu.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10164__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06541_ _02619_ _02827_ _02882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09260_ _04448_ _04583_ _04590_ _01251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06472_ u_cpu.rf_ram.memory\[41\]\[2\] _02840_ _02843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08682__A1 _03703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07485__A2 _03425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05423_ u_cpu.rf_ram.memory\[16\]\[5\] u_cpu.rf_ram.memory\[17\]\[5\] u_cpu.rf_ram.memory\[18\]\[5\]
+ u_cpu.rf_ram.memory\[19\]\[5\] _01508_ _01509_ _02003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__05040__S0 _01529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08211_ u_arbiter.i_wb_cpu_rdt\[18\] _03822_ _03833_ u_arbiter.i_wb_cpu_dbus_dat\[19\]
+ _03861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_60_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09191_ _02768_ _02870_ _04552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05354_ _01463_ _01934_ _01558_ _01935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08142_ _03804_ _03805_ _03809_ _00914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08434__A1 _03701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07237__A2 _03277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05248__A1 _01506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08073_ u_cpu.rf_ram.memory\[122\]\[6\] _03760_ _03767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05285_ u_cpu.rf_ram.memory\[104\]\[3\] u_cpu.rf_ram.memory\[105\]\[3\] u_cpu.rf_ram.memory\[106\]\[3\]
+ u_cpu.rf_ram.memory\[107\]\[3\] _01555_ _01531_ _01867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_119_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07024_ u_cpu.rf_ram.memory\[5\]\[0\] _03167_ _03168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06748__A1 _02885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08975_ u_cpu.rf_ram.memory\[97\]\[4\] _04425_ _04430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05420__A1 _01506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07926_ _03681_ _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09162__A2 _04533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10507__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07857_ _02277_ _03638_ _03640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07173__A1 _02642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06808_ u_cpu.rf_ram.memory\[6\]\[4\] _03039_ _03044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08277__S _02465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05723__A2 _02292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07788_ u_cpu.rf_ram.memory\[36\]\[5\] _03593_ _03599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09527_ _02395_ u_cpu.cpu.genblk3.csr.timer_irq_r _04235_ _04750_ _01358_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_06739_ u_cpu.rf_ram.memory\[77\]\[6\] _02998_ _03005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10657__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09458_ _04628_ _04701_ _04704_ _01335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07476__A2 _03415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08409_ _03910_ _04021_ _04027_ _04028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09389_ u_cpu.rf_ram.memory\[85\]\[4\] _04661_ _04666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05582__S1 _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07228__A2 _03277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05239__A1 _01812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08976__A2 _04425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10302_ _00688_ io_in[4] u_cpu.rf_ram.memory\[12\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08740__S _02335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10037__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10233_ _00619_ io_in[4] u_cpu.rf_ram.memory\[137\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05098__S0 _01576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10164_ _00550_ io_in[4] u_cpu.rf_ram.memory\[72\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07400__A2 _03375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05411__A1 _01465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10095_ _00489_ io_in[4] u_cpu.rf_ram.memory\[53\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10187__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09153__A2 _04523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08900__A2 _04371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05270__S0 _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10997_ _01366_ io_in[4] u_cpu.rf_ram.memory\[27\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05190__A3 _01753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07467__A2 _03415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08664__A1 _03703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05573__S1 _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08416__A1 _03974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07219__A2 _03267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08967__A2 _04425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05559__B _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05070_ _01513_ _01653_ _01654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05089__S0 _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09392__A2 _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05402__A1 _01617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08760_ _02355_ _04296_ _04293_ _04297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05972_ u_cpu.cpu.ctrl.o_ibus_adr\[8\] _02486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09822__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09144__A2 _04523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07711_ _03500_ _03553_ _03556_ _00735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_04923_ _01507_ _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08691_ _04258_ _01014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07155__A1 _03104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09695__A3 u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07642_ u_cpu.rf_ram.memory\[128\]\[4\] _03513_ _03518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04854_ u_cpu.cpu.decode.co_mem_word _01441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05261__S0 _01495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07573_ _03306_ _03475_ _03476_ _00677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09972__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09312_ _04446_ _04613_ _04619_ _01274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06524_ u_cpu.rf_ram.memory\[47\]\[0\] _02872_ _02873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07458__A2 _03405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05469__A1 _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09243_ u_cpu.rf_ram.memory\[106\]\[7\] _04573_ _04581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06455_ u_cpu.rf_ram.memory\[51\]\[3\] _02829_ _02833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05564__S1 _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08407__A1 _03901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05406_ u_cpu.rf_ram.memory\[136\]\[4\] u_cpu.rf_ram.memory\[137\]\[4\] u_cpu.rf_ram.memory\[138\]\[4\]
+ u_cpu.rf_ram.memory\[139\]\[4\] _01634_ _01635_ _01987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09174_ _04542_ _04543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06386_ u_cpu.rf_ram.memory\[42\]\[7\] _02784_ _02792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05337_ _01911_ _01913_ _01915_ _01917_ _01486_ _01918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_08125_ u_cpu.rf_ram.memory\[33\]\[5\] _03790_ _03796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08056_ _03705_ _03750_ _03757_ _00880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05268_ u_cpu.rf_ram.memory\[60\]\[3\] u_cpu.rf_ram.memory\[61\]\[3\] u_cpu.rf_ram.memory\[62\]\[3\]
+ u_cpu.rf_ram.memory\[63\]\[3\] _01496_ _01563_ _01850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07630__A2 _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05188__C _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05641__A1 _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07007_ _03098_ _03157_ _03158_ _00429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05199_ _01775_ _01777_ _01779_ _01781_ _01560_ _01782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_143_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09383__A2 _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08958_ _04413_ _04414_ _04418_ _01121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09135__A2 _04513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07909_ u_cpu.rf_ram.memory\[34\]\[0\] _03672_ _03673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08889_ _02667_ _04361_ _04369_ _01101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_99_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08343__B1 _03958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10920_ _01289_ io_in[4] u_cpu.rf_ram.memory\[59\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07697__A2 _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05252__S0 _01530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10851_ _01220_ io_in[4] u_cpu.rf_ram.memory\[99\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07449__A2 _03405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10782_ _01151_ io_in[4] u_cpu.rf_ram.memory\[96\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05004__S0 _01551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05379__B _01600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05307__S1 _01622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07621__A2 _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08470__S _02466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05632__A1 _01512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09845__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09374__A2 _04651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10216_ _00602_ io_in[4] u_cpu.rf_ram.memory\[138\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07385__A1 _02657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10147_ _00533_ io_in[4] u_cpu.rf_ram.memory\[140\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10822__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05935__A2 _02456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09126__A2 _04513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07137__A1 _03104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10078_ _00472_ io_in[4] u_cpu.rf_ram.memory\[55\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09995__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07688__A2 _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08885__A1 _02657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05699__A1 _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05243__S0 _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10972__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06360__A2 _02770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_63_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08637__A1 _03955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06112__A2 u_arbiter.i_wb_cpu_ibus_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10202__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06240_ _02689_ _02697_ _02703_ _00117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07860__A2 _02309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06171_ _02651_ _02652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05122_ u_cpu.rf_ram.memory\[92\]\[1\] u_cpu.rf_ram.memory\[93\]\[1\] u_cpu.rf_ram.memory\[94\]\[1\]
+ u_cpu.rf_ram.memory\[95\]\[1\] _01562_ _01563_ _01706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_50_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07612__A2 _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10352__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05623__A1 _01548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05053_ _01621_ _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09930_ _00324_ io_in[4] u_cpu.rf_ram.memory\[74\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09365__A2 _04651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09861_ _00255_ io_in[4] u_cpu.rf_ram.memory\[4\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08412__I1 u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06179__A2 _02657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08812_ u_cpu.cpu.ctrl.o_ibus_adr\[14\] _04309_ _04311_ u_cpu.cpu.ctrl.o_ibus_adr\[15\]
+ _04326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_112_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09792_ _00186_ io_in[4] u_cpu.rf_ram.memory\[45\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09117__A2 _04503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08743_ _04284_ _01040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05955_ _02467_ u_cpu.cpu.ctrl.o_ibus_adr\[3\] u_cpu.cpu.ctrl.o_ibus_adr\[2\] _02473_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_39_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05139__B1 _01720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04906_ _01467_ u_cpu.rf_ram_if.wtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__07679__A2 _03533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08674_ _03695_ _04247_ _04249_ _01006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05886_ u_arbiter.i_wb_cpu_rdt\[14\] u_arbiter.i_wb_cpu_dbus_dat\[11\] _02418_ _02429_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_27_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05234__S0 _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07625_ _03506_ _03496_ _03507_ _00698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06351__A2 _02770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08628__A1 _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07556_ u_cpu.rf_ram.memory\[131\]\[1\] _03465_ _03467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06507_ u_cpu.rf_ram.memory\[48\]\[1\] _02861_ _02863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09718__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07487_ _03312_ _03425_ _03428_ _00639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07300__A1 _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09226_ _04450_ _04563_ _04571_ _01236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06438_ u_cpu.rf_ram.memory\[44\]\[5\] _02816_ _02822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07851__A2 _02305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09157_ u_cpu.rf_ram.memory\[104\]\[0\] _04533_ _04534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09053__A1 _04434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06369_ _02781_ _02782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08108_ _03703_ _03780_ _03786_ _00903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09868__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09088_ _04495_ _01174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07603__A2 _03485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05614__A1 _01504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08039_ u_cpu.rf_ram.memory\[11\]\[7\] _03740_ _03748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10845__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11050_ _01419_ io_in[4] u_cpu.rf_ram.memory\[89\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09356__A2 _04641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07367__A1 _03318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10001_ _00395_ io_in[4] u_cpu.rf_ram.memory\[29\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09108__A2 _04503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07119__A1 _03104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10995__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05662__B _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08867__A1 _03703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05225__S0 _01529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10903_ _01272_ io_in[4] u_cpu.rf_ram.memory\[69\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06342__A2 _02756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10225__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10834_ _01203_ io_in[4] u_cpu.rf_ram.memory\[103\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09292__A1 _04444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10765_ _01134_ io_in[4] u_cpu.rf_ram.memory\[94\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08095__A2 _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07842__A2 _03626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10696_ _01066_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10375__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05853__A1 u_arbiter.i_wb_cpu_rdt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09044__A1 _04450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09595__A2 _04782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05605__A1 _01528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09347__A2 _04641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05464__S0 _01496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11000__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06581__A2 _02900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05740_ _01442_ u_arbiter.i_wb_cpu_dbus_dat\[5\] _02314_ u_cpu.cpu.state.init_done
+ _02315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__05216__S0 _01507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05671_ _01465_ _02248_ _02249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_90_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06333__A2 _02756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07410_ u_cpu.rf_ram.memory\[39\]\[0\] _03385_ _03386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11150__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08390_ u_arbiter.i_wb_cpu_rdt\[20\] u_arbiter.i_wb_cpu_rdt\[4\] _02467_ _04010_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_35_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10718__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07341_ _03310_ _03345_ _03347_ _00574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08086__A2 _03770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06097__A1 _02265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07272_ u_cpu.rf_ram.memory\[13\]\[7\] _03297_ _03305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07833__A2 _02780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09011_ u_cpu.rf_ram.memory\[95\]\[0\] _04453_ _04454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06223_ _02666_ _02693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_129_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10868__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06154_ u_cpu.rf_ram.memory\[82\]\[1\] _02628_ _02638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09586__A2 _04782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07597__A1 _02647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05105_ u_cpu.rf_ram.memory\[96\]\[1\] u_cpu.rf_ram.memory\[97\]\[1\] u_cpu.rf_ram.memory\[98\]\[1\]
+ u_cpu.rf_ram.memory\[99\]\[1\] _01567_ _01568_ _01689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08794__B1 _04311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06085_ u_cpu.cpu.ctrl.o_ibus_adr\[29\] u_cpu.cpu.ctrl.o_ibus_adr\[28\] u_cpu.cpu.ctrl.o_ibus_adr\[27\]
+ _02562_ _02577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_105_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09338__A2 _04624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09913_ _00307_ io_in[4] u_cpu.rf_ram.memory\[139\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05036_ _01504_ _01621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_63_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07349__A1 _03318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09844_ _00238_ io_in[4] u_cpu.rf_ram.memory\[47\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08010__A2 _03730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05455__S0 _01551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09775_ _00169_ io_in[4] u_cpu.rf_ram.memory\[42\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_101_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06987_ _03146_ _03147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06572__A2 _02900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10248__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08726_ u_arbiter.i_wb_cpu_dbus_adr\[20\] u_arbiter.i_wb_cpu_dbus_adr\[21\] _02335_
+ _04276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__04877__I _01463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05938_ u_arbiter.i_wb_cpu_ibus_adr\[1\] _02456_ _02459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08849__A1 _02276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08657_ u_cpu.rf_ram.memory\[32\]\[2\] _04237_ _04240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05869_ _02420_ _00094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07521__A1 _03310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06324__A2 _02745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07608_ _03495_ _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08588_ _03908_ _03918_ _04179_ _04180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_41_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10398__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07539_ _03310_ _03455_ _03457_ _00662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_41_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08077__A2 _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09274__A1 _04444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06088__A1 _02397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10550_ _00923_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07824__A2 _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09209_ _02838_ _04349_ _04562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09026__A1 _04450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10481_ _00854_ io_in[4] u_cpu.rf_ram.memory\[121\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09577__A2 _04772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07588__A1 _02731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05657__B _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11102_ _00031_ io_in[0] u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05063__A2 _01647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06260__A1 _02691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09329__A2 _04624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11023__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11033_ _01402_ io_in[4] u_cpu.rf_ram.memory\[98\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08001__A2 _03720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06012__A1 _02456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05446__S0 _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05366__A3 _01927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06315__A2 _02745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10817_ _01186_ io_in[4] u_cpu.rf_ram.memory\[101\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08068__A2 _03760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08312__I0 u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06079__A1 _02402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10748_ _01117_ io_in[4] u_cpu.rf_ram.memory\[93\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07815__A2 _02849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10679_ _01051_ io_in[4] u_cpu.rf_ram.memory\[30\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09568__A2 _04772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07579__A1 _03314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08240__A2 _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06910_ _03098_ _03100_ _03101_ _00389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07890_ _03661_ _03662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06003__A1 _02402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06003__B2 u_arbiter.i_wb_cpu_dbus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05437__S0 _01495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06841_ _02887_ _03059_ _03062_ _00359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07751__A1 _03504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09560_ u_cpu.rf_ram.memory\[26\]\[6\] _04762_ _04769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06772_ _02891_ _03018_ _03023_ _00329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08511_ _03944_ _03975_ _03938_ _04112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05723_ _02295_ _02292_ _02296_ _02298_ _02299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_09491_ u_cpu.cpu.genblk3.csr.mcause3_0\[1\] _04724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10540__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07503__A1 _03310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08442_ _03906_ _03947_ _04051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05654_ u_cpu.rf_ram.memory\[80\]\[7\] u_cpu.rf_ram.memory\[81\]\[7\] u_cpu.rf_ram.memory\[82\]\[7\]
+ u_cpu.rf_ram.memory\[83\]\[7\] _01544_ _01545_ _02232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_23_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09256__A1 _04444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08059__A2 _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08373_ _02466_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[10\] _03995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_51_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05585_ _01638_ _02163_ _01482_ _02164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10690__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07324_ u_cpu.rf_ram.memory\[71\]\[2\] _03335_ _03338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07806__A2 _02927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05817__A1 _01467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09008__A1 _04450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07255_ _03114_ _03287_ _03295_ _00540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06085__A4 _02562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05293__A2 _01874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06206_ u_cpu.rf_ram.memory\[21\]\[1\] _02679_ _02682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06490__A1 _02681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09559__A2 _04762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07186_ u_cpu.rf_ram.memory\[15\]\[0\] _03257_ _03258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11046__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05477__B _01600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06137_ _02606_ u_cpu.rf_ram_if.wen1_r u_cpu.rf_ram_if.rtrig0 u_cpu.rf_ram_if.wen0_r
+ _02622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08231__A2 _03802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05045__A2 _01629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06242__A1 _02691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05676__S0 _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06068_ u_cpu.cpu.ctrl.o_ibus_adr\[26\] _02563_ _02456_ _02564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07990__A1 _03691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06793__A2 _03028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09906__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05019_ _01602_ _01603_ _01604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10070__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05428__S0 _01530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09827_ _00221_ io_in[4] u_cpu.rf_ram.memory\[43\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09758_ _00152_ io_in[4] u_cpu.rf_ram.memory\[80\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08709_ _04267_ _01023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09689_ _04638_ _04832_ _04840_ _01430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08298__A2 _03923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09495__A1 _04723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04859__A2 _01445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10602_ _00975_ io_in[4] u_cpu.cpu.immdec.imm24_20\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05808__A1 _02273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10533_ _00906_ io_in[4] u_cpu.rf_ram.memory\[33\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05284__A2 _01865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06481__A1 _02691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10464_ _00837_ io_in[4] u_cpu.rf_ram.memory\[120\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08222__A2 _03808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10395_ _00768_ io_in[4] u_cpu.rf_ram.memory\[36\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10413__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06784__A2 _03028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11016_ _01385_ io_in[4] u_cpu.rf_ram.memory\[24\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05419__S0 _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10563__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07733__A1 _03504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06536__A2 _02872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09486__A1 _04638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08289__A2 u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09238__A1 _04444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05370_ _01548_ _01950_ _01579_ _01951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11069__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08461__A2 _04068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05275__A2 _01856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07040_ _02780_ _02827_ _03176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09929__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10093__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09410__A1 _04634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08213__A2 _03808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08991_ _02641_ _04440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06775__A2 _03018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07972__A1 _03691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10906__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07942_ _03510_ _03682_ _03690_ _00833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07873_ u_cpu.rf_ram.memory\[92\]\[0\] _03652_ _03653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06527__A2 _02872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09612_ u_cpu.rf_ram.memory\[0\]\[5\] _04792_ _04798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_95_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06824_ u_cpu.rf_ram.memory\[68\]\[3\] _03049_ _03053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09543_ _04636_ _04752_ _04759_ _01365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06755_ u_cpu.rf_ram.memory\[74\]\[5\] _03008_ _03014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05706_ _01441_ u_cpu.cpu.bne_or_bge _02282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09474_ _04626_ _04711_ _04713_ _01342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06686_ u_cpu.rf_ram.memory\[119\]\[7\] _02967_ _02975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08425_ u_cpu.rf_ram.memory\[114\]\[0\] _04041_ _04042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05637_ u_cpu.rf_ram.memory\[104\]\[7\] u_cpu.rf_ram.memory\[105\]\[7\] u_cpu.rf_ram.memory\[106\]\[7\]
+ u_cpu.rf_ram.memory\[107\]\[7\] _01555_ _01531_ _02215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_12_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08356_ _03914_ _03908_ _03912_ _03980_ _03896_ _03981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__06147__I _02631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05568_ u_cpu.rf_ram.memory\[84\]\[6\] u_cpu.rf_ram.memory\[85\]\[6\] u_cpu.rf_ram.memory\[86\]\[6\]
+ u_cpu.rf_ram.memory\[87\]\[6\] _01507_ _01605_ _02147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_138_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07307_ _03312_ _03325_ _03328_ _00559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08287_ _03914_ _03903_ _03915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05499_ _01465_ _02078_ _02079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_137_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10436__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07238_ _02814_ _02976_ _03286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07169_ _02632_ _03247_ _03248_ _00501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08204__A2 _03835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10180_ _00566_ io_in[4] u_cpu.rf_ram.memory\[71\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10586__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06766__A2 _03018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08507__A3 _04093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07715__A1 _03504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06518__A2 _02861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08738__S _02335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07191__A2 _03257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09468__A1 _04638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08140__A1 _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08443__A2 _04051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05257__A2 _01838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06454__A1 _02683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10516_ _00889_ io_in[4] u_cpu.rf_ram.memory\[122\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10929__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10447_ _00820_ io_in[4] u_cpu.rf_ram.memory\[34\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10378_ _00751_ io_in[4] u_cpu.rf_ram.memory\[38\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06757__A2 _03008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06509__A2 _02861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05980__A3 _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04870_ _01444_ _01445_ _01457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07182__A2 _03247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10309__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06540_ _02631_ _02881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__04975__I _01540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08131__A1 u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06471_ _02681_ _02840_ _02842_ _00209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08682__A2 _04247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10459__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08210_ u_arbiter.i_wb_cpu_dbus_dat\[18\] _03835_ _03860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05422_ _01513_ _02001_ _02002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05040__S1 _01500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09190_ _04450_ _04543_ _04551_ _01220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_18_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08141_ u_arbiter.i_wb_cpu_rdt\[0\] _03807_ _03808_ u_arbiter.i_wb_cpu_dbus_dat\[0\]
+ _03809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_53_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05353_ u_cpu.rf_ram.memory\[44\]\[4\] u_cpu.rf_ram.memory\[45\]\[4\] u_cpu.rf_ram.memory\[46\]\[4\]
+ u_cpu.rf_ram.memory\[47\]\[4\] _01555_ _01531_ _01934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09751__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09631__A1 _04634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08434__A2 _04041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05248__A2 _01829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06445__A1 _02728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08072_ _03703_ _03760_ _03766_ _00887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05284_ _01512_ _01865_ _01866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06996__A2 _03147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07023_ _03166_ _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_115_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06748__A2 _03008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05755__B u_arbiter.i_wb_cpu_ibus_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08974_ _03699_ _04425_ _04429_ _01126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08131__B _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07925_ _02675_ _02965_ _03681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05420__A2 _01999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07856_ u_cpu.cpu.alu.i_rs1 _03638_ _03639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07173__A2 _03247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08370__A1 _03956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06807_ _02647_ _03039_ _03043_ _00344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_83_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07787_ _03504_ _03593_ _03598_ _00769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06586__B _02910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04999_ _01492_ _01521_ _01542_ _01583_ _01584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_45_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05490__B _01481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09526_ u_cpu.cpu.genblk3.csr.o_new_irq _03611_ _04750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06738_ _02893_ _02998_ _03004_ _00314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08122__A1 _03699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09457_ u_cpu.rf_ram.memory\[87\]\[2\] _04701_ _04704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06669_ _02728_ _02624_ _02729_ _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__08673__A2 _04247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08408_ _03938_ _04023_ _04026_ _03944_ _04027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_61_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09388_ _04630_ _04661_ _04665_ _01304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08339_ _03964_ _03965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08425__A2 _04041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05239__A2 _01821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10301_ _00687_ io_in[4] u_cpu.rf_ram.memory\[12\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04998__A1 _01490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10232_ _00618_ io_in[4] u_cpu.rf_ram.memory\[137\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06739__A2 _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07936__A1 _03504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05098__S1 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10163_ _00549_ io_in[4] u_cpu.rf_ram.memory\[72\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05411__A2 _01991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05384__C _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09689__A1 _04638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10094_ _00488_ io_in[4] u_cpu.rf_ram.memory\[53\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08361__A1 _03915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07164__A2 _03237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05270__S1 _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10601__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10996_ _01365_ io_in[4] u_cpu.rf_ram.memory\[27\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08113__A1 _02695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09774__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06124__B1 _02608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08664__A2 _04237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06675__A1 _02885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10751__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09613__A1 _02689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06978__A2 _03137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11107__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05089__S1 _01531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05402__A2 _01982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05971_ _02456_ _02484_ _02485_ _00065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10131__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07710_ u_cpu.rf_ram.memory\[124\]\[2\] _03553_ _03556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04922_ _01494_ _01507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_38_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08690_ u_arbiter.i_wb_cpu_dbus_adr\[2\] u_arbiter.i_wb_cpu_dbus_adr\[3\] _04257_
+ _04258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08378__S _02466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07155__A2 _03237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07641_ _03502_ _03513_ _03517_ _00704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04853_ u_cpu.cpu.immdec.imm24_20\[0\] _01440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_93_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06902__A2 _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10281__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05261__S1 _01499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07572_ u_cpu.rf_ram.memory\[130\]\[0\] _03475_ _03476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08104__A1 _03699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09311_ u_cpu.rf_ram.memory\[69\]\[5\] _04613_ _04619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06523_ _02871_ _02872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_62_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08655__A2 _04237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09242_ _04448_ _04573_ _04580_ _01243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05469__A2 _02048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06666__A1 _02895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06454_ _02683_ _02829_ _02832_ _00202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05405_ _01966_ _01985_ _01471_ _01986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09173_ _02825_ _04349_ _04542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08407__A2 _03975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06385_ _02691_ _02784_ _02791_ _00174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06418__A1 _02687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08124_ _03701_ _03790_ _03795_ _00910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05336_ _01506_ _01916_ _01519_ _01917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_135_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08055_ u_cpu.rf_ram.memory\[112\]\[6\] _03750_ _03757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07091__A1 _03112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05267_ _01842_ _01844_ _01846_ _01848_ _01560_ _01849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_134_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07006_ u_cpu.rf_ram.memory\[19\]\[0\] _03157_ _03158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05641__A2 _02218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05198_ _01566_ _01780_ _01558_ _01781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07918__A1 _03504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08591__A1 _03947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07394__A2 _03375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08957_ _03956_ _04417_ _04418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07908_ _03671_ _03672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10624__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08888_ u_cpu.rf_ram.memory\[3\]\[7\] _04361_ _04369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08343__A1 _02313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07146__A2 _03227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08343__B2 _03959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07839_ u_cpu.rf_ram.memory\[90\]\[2\] _03626_ _03629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09797__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08894__A2 _04371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10850_ _01219_ io_in[4] u_cpu.rf_ram.memory\[99\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05252__S1 _01532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04904__A1 _01473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09509_ _04736_ u_cpu.cpu.genblk3.csr.mcause31 _04737_ _04738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10781_ _01150_ io_in[4] u_cpu.rf_ram.memory\[96\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10774__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05004__S1 _01524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10004__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10154__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10215_ _00601_ io_in[4] u_cpu.rf_ram.memory\[138\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07385__A2 _03365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10146_ _00532_ io_in[4] u_cpu.rf_ram.memory\[141\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05396__A1 _01621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10077_ _00471_ io_in[4] u_cpu.rf_ram.memory\[55\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08334__A1 _03936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07137__A2 _03227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08885__A2 _04361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05243__S1 _01509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05699__A2 _02274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10979_ _01348_ io_in[4] u_cpu.rf_ram.memory\[88\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06170_ _02650_ _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09062__A2 _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05121_ _01490_ _01695_ _01704_ _01705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__07073__A1 _03112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05052_ _01465_ _01636_ _01637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_125_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09860_ _00254_ io_in[4] u_cpu.rf_ram.memory\[4\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10647__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07376__A2 _03365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08811_ _04325_ _01067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__05387__A1 _01464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09791_ _00185_ io_in[4] u_cpu.rf_ram.memory\[45\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08742_ u_arbiter.i_wb_cpu_dbus_adr\[28\] u_arbiter.i_wb_cpu_dbus_adr\[29\] _02335_
+ _04284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05954_ _02456_ _02471_ _02472_ _00061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09505__B _04723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08325__A1 _02265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07128__A2 _03217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04905_ _01465_ _01491_ _00025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_61_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08673_ u_cpu.rf_ram.memory\[31\]\[1\] _04247_ _04249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10797__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05885_ _02428_ _00033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08876__A2 _04361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07624_ u_cpu.rf_ram.memory\[22\]\[5\] _03496_ _03507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06887__A1 _02897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05234__S1 _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07555_ _03306_ _03465_ _03466_ _00669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08628__A2 _02414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10027__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04993__S0 _01576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06639__A1 _02887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06506_ _02669_ _02861_ _02862_ _00224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07486_ u_cpu.rf_ram.memory\[135\]\[2\] _03425_ _03428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07300__A2 _02838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09225_ u_cpu.rf_ram.memory\[105\]\[7\] _04563_ _04571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06437_ _02687_ _02816_ _02821_ _00196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09156_ _04532_ _04533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05199__C _01560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06368_ u_cpu.cpu.immdec.imm11_7\[2\] u_cpu.cpu.immdec.imm11_7\[4\] _02622_ _02729_
+ _02781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__09053__A2 _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10177__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08107_ u_cpu.rf_ram.memory\[116\]\[5\] _03780_ _03786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05319_ _01465_ _01900_ _01901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09087_ u_arbiter.i_wb_cpu_rdt\[25\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[9\]
+ _04485_ _04495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08800__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06299_ u_cpu.rf_ram.memory\[1\]\[5\] _02733_ _02739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06811__A1 _02657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08038_ _02662_ _03740_ _03747_ _00872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05614__A2 _02191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10000_ _00394_ io_in[4] u_cpu.rf_ram.memory\[29\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08564__A1 _02392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07367__A2 _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09989_ _00383_ io_in[4] u_cpu.rf_ram.memory\[64\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08316__A1 _02465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07119__A2 _03217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08867__A2 _04351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05225__S1 _01500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10902_ _01271_ io_in[4] u_cpu.rf_ram.memory\[69\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08746__S _02335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10833_ _01202_ io_in[4] u_cpu.rf_ram.memory\[103\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05550__A1 _01566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08619__A2 _03955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04984__S0 _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10764_ _01133_ io_in[4] u_cpu.rf_ram.memory\[94\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09292__A2 _04603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10695_ _01065_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05853__A2 _02389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09812__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09044__A2 _04463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07055__A1 _03112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09962__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08555__A1 _03935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07358__A2 _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06030__A2 _02397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10129_ _00006_ io_in[4] u_cpu.rf_ram.rdata\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05464__S1 _01594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08307__A1 _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08858__A2 _04351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05216__S1 _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06869__A1 _02897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05670_ u_cpu.rf_ram.memory\[128\]\[7\] u_cpu.rf_ram.memory\[129\]\[7\] u_cpu.rf_ram.memory\[130\]\[7\]
+ u_cpu.rf_ram.memory\[131\]\[7\] _01641_ _01642_ _02248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_17_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07530__A2 _03445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05541__A1 _01490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07340_ u_cpu.rf_ram.memory\[70\]\[1\] _03345_ _03347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__04983__I _01498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09283__A2 _04603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07271_ _02662_ _03297_ _03304_ _00547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09010_ _04452_ _04453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06222_ _02691_ _02679_ _02692_ _00110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09035__A2 _04463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06153_ _02636_ _02637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05104_ _01571_ _01687_ _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07597__A2 _03485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06084_ _02389_ u_scanchain_local.module_data_in\[67\] _02576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05035_ _01612_ _01614_ _01616_ _01619_ _01486_ _01620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_99_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09912_ _00306_ io_in[4] u_cpu.rf_ram.memory\[139\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08546__A1 _01444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07349__A2 _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09843_ _00237_ io_in[4] u_cpu.rf_ram.memory\[47\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05455__S1 _01524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09774_ _00168_ io_in[4] u_cpu.rf_ram.memory\[42\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06986_ _02814_ _02827_ _03146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05482__C _01486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05937_ _02403_ u_scanchain_local.module_data_in\[38\] _02458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08725_ _04275_ _01031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08849__A2 _02334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08656_ _03695_ _04237_ _04239_ _00998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05868_ u_arbiter.i_wb_cpu_rdt\[5\] u_arbiter.i_wb_cpu_dbus_dat\[2\] _02418_ _02420_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__05907__I0 u_arbiter.i_wb_cpu_rdt\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07521__A2 _03445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07607_ _02677_ _03037_ _03495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08587_ _03924_ _04052_ _03915_ _04179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05799_ _02273_ u_cpu.rf_ram.rdata\[2\] _02371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07538_ u_cpu.rf_ram.memory\[132\]\[1\] _03455_ _03457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09835__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09274__A2 _04593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07469_ _03312_ _03415_ _03418_ _00631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05003__B _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09208_ _04450_ _04553_ _04561_ _01228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10812__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10480_ _00853_ io_in[4] u_cpu.rf_ram.memory\[121\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09026__A2 _04453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09139_ u_cpu.rf_ram.memory\[103\]\[0\] _04523_ _04524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07037__A1 _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09985__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08234__B1 _03874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07588__A2 _02814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11101_ _00030_ io_in[0] u_arbiter.i_wb_cpu_rdt\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10962__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06260__A2 _02707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11032_ _01401_ io_in[4] u_cpu.rf_ram.memory\[98\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05673__B _01482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05446__S1 _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07760__A2 _03583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05771__A1 u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07512__A2 _03435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10342__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10816_ _01185_ io_in[4] u_cpu.rf_ram.memory\[101\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09265__A2 _04593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10747_ _01116_ io_in[4] u_cpu.rf_ram.memory\[93\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10492__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05826__A2 _01467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09017__A2 _04453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10678_ _01050_ io_in[4] u_cpu.rf_ram.memory\[30\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05382__S0 _01576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07579__A2 _03475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06251__A2 _02707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08528__A1 _03923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09708__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06840_ u_cpu.rf_ram.memory\[67\]\[2\] _03059_ _03062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__04978__I _01499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05437__S1 _01499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07751__A2 _03573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06771_ u_cpu.rf_ram.memory\[76\]\[4\] _03018_ _03023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05762__A1 _02322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08510_ _03932_ _03988_ _04111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05722_ _02259_ _02297_ _02298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09490_ _04722_ _04723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_63_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09858__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07503__A2 _03435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08441_ u_arbiter.i_wb_cpu_rdt\[26\] u_arbiter.i_wb_cpu_rdt\[10\] _02466_ _04050_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05653_ _01597_ _02230_ _01600_ _02231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_63_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09502__C _02305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04948__S0 _01530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08372_ _03965_ _03961_ _03994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10835__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05584_ u_cpu.rf_ram.memory\[132\]\[6\] u_cpu.rf_ram.memory\[133\]\[6\] u_cpu.rf_ram.memory\[134\]\[6\]
+ u_cpu.rf_ram.memory\[135\]\[6\] _01634_ _01635_ _02163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09256__A2 _04583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07323_ _03310_ _03335_ _03337_ _00566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07267__A1 _02652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07254_ u_cpu.rf_ram.memory\[140\]\[7\] _03287_ _03295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05817__A2 _02369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05373__S0 _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09008__A2 _04436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06205_ _02636_ _02681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07019__A1 _03112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10985__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07185_ _03256_ _03257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06490__A2 _02851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08767__A1 _03695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06136_ u_cpu.cpu.immdec.imm11_7\[4\] _02621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06242__A2 _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06067_ _02561_ _02554_ _02563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05676__S1 _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10215__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08519__A1 _03958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05049__I _01522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07990__A2 _03720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05018_ u_cpu.rf_ram.memory\[112\]\[0\] u_cpu.rf_ram.memory\[113\]\[0\] u_cpu.rf_ram.memory\[114\]\[0\]
+ u_cpu.rf_ram.memory\[115\]\[0\] _01544_ _01545_ _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_132_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05493__B _01471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09826_ _00220_ io_in[4] u_cpu.rf_ram.memory\[43\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05428__S1 _01532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07742__A2 _03573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10365__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09757_ _00151_ io_in[4] u_cpu.rf_ram.memory\[7\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06969_ _03136_ _03137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_104_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08708_ u_arbiter.i_wb_cpu_dbus_adr\[11\] u_arbiter.i_wb_cpu_dbus_adr\[12\] _04257_
+ _04267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08296__S _02464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09688_ u_cpu.rf_ram.memory\[23\]\[7\] _04832_ _04840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08298__A3 _03924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08639_ _02305_ _01440_ _03896_ _04227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09247__A2 _04583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10601_ _00974_ io_in[4] u_cpu.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10532_ _00905_ io_in[4] u_cpu.rf_ram.memory\[116\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10463_ _00836_ io_in[4] u_cpu.rf_ram.memory\[120\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06481__A2 _02840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08758__A1 u_arbiter.i_wb_cpu_dbus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05116__S0 _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10394_ _00767_ io_in[4] u_cpu.rf_ram.memory\[36\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06233__A2 _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11140__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07981__A2 _03710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10708__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11015_ _01384_ io_in[4] u_cpu.rf_ram.memory\[24\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05419__S1 _01509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07733__A2 _03563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08930__A1 _03932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05744__A1 _01445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10858__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09486__A2 _04711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07497__A1 _03322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09238__A2 _04573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07249__A1 _03108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08297__I0 u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05578__B _01600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06472__A2 _02840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10238__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05107__S0 _01551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09410__A2 _04671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06224__A2 _02679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07421__A1 _03318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08990_ _04438_ _04436_ _04439_ _01132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07972__A2 _03710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07941_ u_cpu.rf_ram.memory\[117\]\[7\] _03682_ _03690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10388__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07872_ _03651_ _03652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08921__A1 _03703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07724__A2 _03563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09611_ _02687_ _04792_ _04797_ _01395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06823_ _02887_ _03049_ _03052_ _00351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05735__A1 _02285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09542_ u_cpu.rf_ram.memory\[27\]\[6\] _04752_ _04759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06754_ _02891_ _03008_ _03013_ _00321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09477__A2 _04711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05705_ _02259_ _02261_ _02281_ _00021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06685_ _02895_ _02967_ _02974_ _00291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09473_ u_cpu.rf_ram.memory\[88\]\[1\] _04711_ _04713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05636_ _01512_ _02213_ _02214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08424_ _04040_ _04041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09229__A2 _04573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11013__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08355_ _02909_ u_arbiter.i_wb_cpu_rdt\[5\] _03979_ _03980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_11_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05567_ _01602_ _02145_ _02146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07306_ u_cpu.rf_ram.memory\[73\]\[2\] _03325_ _03328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08286_ _02909_ u_arbiter.i_wb_cpu_rdt\[0\] _03913_ _03914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05498_ u_cpu.rf_ram.memory\[128\]\[5\] u_cpu.rf_ram.memory\[129\]\[5\] u_cpu.rf_ram.memory\[130\]\[5\]
+ u_cpu.rf_ram.memory\[131\]\[5\] _01641_ _01642_ _02078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07237_ _03114_ _03277_ _03285_ _00532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06463__A2 _02829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07168_ u_cpu.rf_ram.memory\[9\]\[0\] _03247_ _03248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09401__A2 _04671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06215__A2 _02679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06119_ u_cpu.cpu.immdec.imm11_7\[4\] _02603_ _02604_ _02598_ _02605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_133_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07099_ _03102_ _03207_ _03209_ _00470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07715__A2 _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09809_ _00203_ io_in[4] u_cpu.rf_ram.memory\[51\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05726__A1 _01460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09468__A2 _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07479__A1 _03322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08140__A2 _03802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06151__A1 _02611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09640__A2 _04812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10515_ _00888_ io_in[4] u_cpu.rf_ram.memory\[122\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05398__B _01519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06454__A2 _02829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10446_ _00819_ io_in[4] u_cpu.rf_ram.memory\[34\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10530__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06206__A2 _02679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07403__A1 _03318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10377_ _00750_ io_in[4] u_cpu.rf_ram.memory\[38\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10680__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07706__A2 _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08903__A1 _02657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05717__A1 u_cpu.cpu.decode.op26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09459__A2 _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11036__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08131__A2 _02355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06470_ u_cpu.rf_ram.memory\[41\]\[1\] _02840_ _02842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06142__A1 _02619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05421_ u_cpu.rf_ram.memory\[20\]\[5\] u_cpu.rf_ram.memory\[21\]\[5\] u_cpu.rf_ram.memory\[22\]\[5\]
+ u_cpu.rf_ram.memory\[23\]\[5\] _01497_ _01501_ _02001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_18_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06693__A2 _02978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10060__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08140_ _03807_ _03802_ _03808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__04991__I _01495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05352_ _01505_ _01932_ _01933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09631__A2 _04802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08071_ u_cpu.rf_ram.memory\[122\]\[5\] _03760_ _03766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06445__A2 u_cpu.cpu.immdec.imm11_7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07642__A1 u_cpu.rf_ram.memory\[128\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05283_ u_cpu.rf_ram.memory\[108\]\[3\] u_cpu.rf_ram.memory\[109\]\[3\] u_cpu.rf_ram.memory\[110\]\[3\]
+ u_cpu.rf_ram.memory\[111\]\[3\] _01529_ _01500_ _01865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08690__I0 u_arbiter.i_wb_cpu_dbus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07022_ _02675_ _02731_ _03166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08198__A2 _03835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09508__B _02303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08973_ u_cpu.rf_ram.memory\[97\]\[3\] _04425_ _04429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05500__S0 _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08131__C _02291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07924_ _03510_ _03672_ _03680_ _00825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07855_ u_cpu.cpu.bne_or_bge _01442_ _01441_ _03638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05708__A1 _01442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06806_ u_cpu.rf_ram.memory\[6\]\[3\] _03039_ _03043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05771__B _01442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06381__A1 _02687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04998_ _01490_ _01561_ _01582_ _01583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_71_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07786_ u_cpu.rf_ram.memory\[36\]\[4\] _03593_ _03598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09525_ _03966_ _04749_ _01357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06737_ u_cpu.rf_ram.memory\[77\]\[5\] _02998_ _03004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08122__A2 _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10403__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09456_ _04626_ _04701_ _04703_ _01334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06133__A1 _01500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06668_ _02897_ _02956_ _02964_ _00284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08407_ _03901_ _03975_ _04025_ _04026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05619_ _02190_ _02192_ _02194_ _02196_ _01560_ _02197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__06684__A2 _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09387_ u_cpu.rf_ram.memory\[85\]\[3\] _04661_ _04665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06599_ _01441_ _02309_ _02922_ _02923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_138_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08338_ _03904_ _03911_ _03964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_137_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09622__A2 _04802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10553__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06436__A2 _02816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08269_ _03896_ _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08830__B1 _04329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06107__B _02596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10300_ _00686_ io_in[4] u_cpu.rf_ram.memory\[12\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_4_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04998__A2 _01561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09386__A1 _04628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08189__A2 _03835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10231_ _00617_ io_in[4] u_cpu.rf_ram.memory\[137\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07936__A2 _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10162_ _00548_ io_in[4] u_cpu.rf_ram.memory\[13\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10093_ _00487_ io_in[4] u_cpu.rf_ram.memory\[53\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09689__A2 _04832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11059__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08361__A2 _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10995_ _01364_ io_in[4] u_cpu.rf_ram.memory\[27\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09919__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10083__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08113__A2 _02782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09310__A1 _04444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08484__S _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06124__A1 _02606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05558__S0 _01576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06124__B2 _02264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05901__S _02431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06675__A2 _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08416__A3 _04024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09613__A2 _04792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07624__A1 u_cpu.rf_ram.memory\[22\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10429_ _00802_ io_in[4] u_cpu.rf_ram.memory\[92\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07927__A2 _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05938__A1 u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05970_ _02418_ u_scanchain_local.module_data_in\[44\] _02398_ u_arbiter.i_wb_cpu_dbus_adr\[7\]
+ _02485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_39_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_04921_ _01505_ _01506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10426__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04852_ u_cpu.cpu.csr_imm _01439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__04986__I _01463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07640_ u_cpu.rf_ram.memory\[128\]\[3\] _03513_ _03517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06363__A1 _02691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05410__I0 u_cpu.rf_ram.memory\[128\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07571_ _03474_ _03475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08104__A2 _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06522_ _02782_ _02870_ _02871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09310_ _04444_ _04613_ _04618_ _01273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05549__S0 _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10576__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09241_ u_cpu.rf_ram.memory\[106\]\[6\] _04573_ _04580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06453_ u_cpu.rf_ram.memory\[51\]\[2\] _02829_ _02832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06666__A2 _02956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04935__B _01519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05404_ _01492_ _01975_ _01984_ _01985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09172_ _04450_ _04533_ _04541_ _01212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06384_ u_cpu.rf_ram.memory\[42\]\[6\] _02784_ _02791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09604__A2 _04792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08123_ u_cpu.rf_ram.memory\[33\]\[4\] _03790_ _03795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05335_ u_cpu.rf_ram.memory\[16\]\[4\] u_cpu.rf_ram.memory\[17\]\[4\] u_cpu.rf_ram.memory\[18\]\[4\]
+ u_cpu.rf_ram.memory\[19\]\[4\] _01508_ _01509_ _01916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06418__A2 _02805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08812__B1 _04311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08054_ _03703_ _03750_ _03756_ _00879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05266_ _01554_ _01847_ _01558_ _01848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07091__A2 _03197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07005_ _03156_ _03157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09368__A1 _02642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05197_ u_cpu.rf_ram.memory\[104\]\[2\] u_cpu.rf_ram.memory\[105\]\[2\] u_cpu.rf_ram.memory\[106\]\[2\]
+ u_cpu.rf_ram.memory\[107\]\[2\] _01555_ _01531_ _01780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_1_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07918__A2 _03672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08040__A1 _02667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08591__A2 _03904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08956_ _03947_ _04031_ _03969_ _03970_ _04416_ _04417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_88_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05057__I _01622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07907_ _02619_ _02782_ _03671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08887_ _02662_ _04361_ _04368_ _01100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_57_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08343__A2 _03956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07838_ _03498_ _03626_ _03628_ _00790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10919__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04904__A2 _01482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07769_ _03504_ _03583_ _03588_ _00761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09508_ _02263_ _02297_ _02303_ _04737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10780_ _01149_ io_in[4] u_cpu.rf_ram.memory\[96\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09439_ u_cpu.rf_ram.memory\[111\]\[2\] _04691_ _04694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06657__A2 _02956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06409__A2 _02805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07082__A2 _03197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05093__A1 _01464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07909__A2 _03672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10214_ _00600_ io_in[4] u_cpu.rf_ram.memory\[138\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06042__B1 _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10145_ _00531_ io_in[4] u_cpu.rf_ram.memory\[141\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10449__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06593__A1 u_arbiter.i_wb_cpu_dbus_dat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05396__A2 _01976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10076_ _00470_ io_in[4] u_cpu.rf_ram.memory\[55\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09531__A1 _04622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09741__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08334__A2 _03938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10599__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06896__A2 _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08098__A1 _03691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09891__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10978_ _01347_ io_in[4] u_cpu.rf_ram.memory\[88\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06648__A2 _02945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05120_ _01697_ _01699_ _01701_ _01703_ _01581_ _01704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_7_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08270__A1 _02465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07073__A2 _03187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05084__A1 _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05051_ u_cpu.rf_ram.memory\[136\]\[0\] u_cpu.rf_ram.memory\[137\]\[0\] u_cpu.rf_ram.memory\[138\]\[0\]
+ u_cpu.rf_ram.memory\[139\]\[0\] _01634_ _01635_ _01636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06820__A2 _03049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08022__A1 _02667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08810_ u_cpu.cpu.ctrl.o_ibus_adr\[13\] _04309_ _04311_ u_cpu.cpu.ctrl.o_ibus_adr\[14\]
+ _04325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08573__A2 _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09790_ _00184_ io_in[4] u_cpu.rf_ram.memory\[45\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05387__A2 _01967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08741_ _04283_ _01039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05953_ _02389_ u_scanchain_local.module_data_in\[40\] _02398_ u_arbiter.i_wb_cpu_dbus_adr\[3\]
+ _02472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__08325__A2 _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09522__A1 u_cpu.cpu.genblk3.csr.mstatus_mie vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_04904_ _01473_ _01482_ _01486_ _01490_ _01491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_94_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08672_ _03691_ _04247_ _04248_ _01005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05884_ u_arbiter.i_wb_cpu_rdt\[13\] u_arbiter.i_wb_cpu_dbus_dat\[10\] _02418_ _02428_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06187__I1 _02368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07623_ _02656_ _03506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06887__A2 _03079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07554_ u_cpu.rf_ram.memory\[131\]\[0\] _03465_ _03466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04993__S1 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06505_ u_cpu.rf_ram.memory\[48\]\[0\] _02861_ _02862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07836__A1 _03494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06639__A2 _02945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07485_ _03310_ _03425_ _03427_ _00638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08137__B _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09224_ _04448_ _04563_ _04570_ _01235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06436_ u_cpu.rf_ram.memory\[44\]\[4\] _02816_ _02821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09589__A1 _04628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09155_ _02954_ _04349_ _04532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06367_ _02618_ _02779_ _02780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08106_ _03701_ _03780_ _03785_ _00902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05318_ u_cpu.rf_ram.memory\[128\]\[3\] u_cpu.rf_ram.memory\[129\]\[3\] u_cpu.rf_ram.memory\[130\]\[3\]
+ u_cpu.rf_ram.memory\[131\]\[3\] _01634_ _01635_ _01900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_135_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08261__A1 _03703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07064__A2 _03187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09086_ _04494_ _01173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06298_ _02652_ _02733_ _02738_ _00140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05075__A1 _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05249_ _01824_ _01826_ _01828_ _01830_ _01486_ _01831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_08037_ u_cpu.rf_ram.memory\[11\]\[6\] _03740_ _03747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06811__A2 _03039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05870__I0 u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06171__I _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08564__A2 _02320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09764__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09988_ _00382_ io_in[4] u_cpu.rf_ram.memory\[64\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06575__A1 _02647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08939_ _03932_ _04009_ _04401_ _03897_ _04402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10741__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08316__A2 _02416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06120__B _02392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10901_ _01270_ io_in[4] u_cpu.rf_ram.memory\[69\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06878__A2 _03079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04889__A1 u_cpu.cpu.decode.op26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10832_ _01201_ io_in[4] u_cpu.rf_ram.memory\[103\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10891__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04984__S1 _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10763_ _01132_ io_in[4] u_cpu.rf_ram.memory\[94\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10694_ _01064_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10121__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07055__A2 _03177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05066__A1 _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06802__A2 _03039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10271__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08004__A1 _03707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08555__A2 _03962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06566__A1 _02717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10128_ _00005_ io_in[4] u_cpu.rf_ram.rdata\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08307__A2 u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10059_ _00453_ io_in[4] u_cpu.rf_ram.memory\[57\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06318__A1 _02652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06869__A2 _03069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05541__A2 _02110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07818__A1 _03494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07270_ u_cpu.rf_ram.memory\[13\]\[6\] _03297_ _03304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08491__A1 _03963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06221_ u_cpu.rf_ram.memory\[21\]\[6\] _02679_ _02692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10614__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06152_ _02635_ _02636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07046__A2 _03177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05103_ u_cpu.rf_ram.memory\[100\]\[1\] u_cpu.rf_ram.memory\[101\]\[1\] u_cpu.rf_ram.memory\[102\]\[1\]
+ u_cpu.rf_ram.memory\[103\]\[1\] _01572_ _01573_ _01687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09787__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08794__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06083_ _02463_ _02574_ _02575_ _00089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05034_ _01617_ _01618_ _01607_ _01619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09911_ _00305_ io_in[4] u_cpu.rf_ram.memory\[139\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10764__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08546__A2 _02265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09842_ _00236_ io_in[4] u_cpu.rf_ram.memory\[47\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09773_ _00167_ io_in[4] u_cpu.rf_ram.memory\[78\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06985_ _03114_ _03137_ _03145_ _00420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08724_ u_arbiter.i_wb_cpu_dbus_adr\[19\] u_arbiter.i_wb_cpu_dbus_adr\[20\] _02335_
+ _04275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_37_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05936_ _02454_ _02457_ _00057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08655_ u_cpu.rf_ram.memory\[32\]\[1\] _04237_ _04239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05867_ _02419_ _00093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_81_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05907__I1 u_arbiter.i_wb_cpu_dbus_dat\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07606_ _02631_ _03494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08586_ _03986_ _03906_ _04177_ _04178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_81_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05798_ _02272_ _02369_ _02370_ _00015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_53_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10144__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07537_ _03306_ _03455_ _03456_ _00661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07809__A1 _02395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07468_ u_cpu.rf_ram.memory\[136\]\[2\] _03415_ _03418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09207_ u_cpu.rf_ram.memory\[79\]\[7\] _04553_ _04561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06419_ u_cpu.rf_ram.memory\[45\]\[5\] _02805_ _02811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07399_ _03314_ _03375_ _03379_ _00600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10294__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09138_ _04522_ _04523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07037__A2 _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08234__A1 u_arbiter.i_wb_cpu_rdt\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05048__A1 _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09069_ u_arbiter.i_wb_cpu_rdt\[16\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[0\]
+ _04485_ _04486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06796__A1 _02897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06115__B _02599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11100_ _00029_ io_in[0] u_arbiter.i_wb_cpu_rdt\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11031_ _01400_ io_in[4] u_cpu.rf_ram.memory\[98\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05220__A1 _01621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05771__A2 _02277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06720__A1 _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10815_ _01184_ io_in[4] u_cpu.rf_ram.memory\[101\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08848__I0 _02363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10637__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10746_ _01115_ io_in[4] u_cpu.rf_ram.memory\[93\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08473__A1 _03941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10677_ _01049_ io_in[4] u_cpu.rf_ram.memory\[30\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05382__S1 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07028__A2 _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05039__A1 _01621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10787__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08776__A2 _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08528__A2 _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10017__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06539__A1 _02693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07200__A2 _03257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05211__A1 _01464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06770_ _02889_ _03018_ _03022_ _00328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10167__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05721_ _01448_ u_cpu.cpu.decode.co_ebreak _01447_ _02297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_64_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08440_ _03707_ _04041_ _04049_ _00972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04994__I _01518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05652_ u_cpu.rf_ram.memory\[88\]\[7\] u_cpu.rf_ram.memory\[89\]\[7\] u_cpu.rf_ram.memory\[90\]\[7\]
+ u_cpu.rf_ram.memory\[91\]\[7\] _01598_ _01556_ _02230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_36_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06187__S _02611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06711__A1 u_cpu.rf_ram.memory\[139\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04948__S1 _01532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08371_ _02286_ _03956_ _03993_ _00959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05583_ _01465_ _02161_ _02162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_32_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07322_ u_cpu.rf_ram.memory\[71\]\[1\] _03335_ _03337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07267__A2 _03297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08464__A1 _04019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05278__A1 _01492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07253_ _03112_ _03287_ _03294_ _00539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05373__S1 _01531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06204_ _02669_ _02679_ _02680_ _00104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07184_ _02731_ _02870_ _03256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07019__A2 _03157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08767__A2 _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06135_ u_cpu.cpu.immdec.imm11_7\[2\] _02608_ _02620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06778__A1 _02897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06066_ _02560_ _02561_ _02555_ _02548_ _02562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__08519__A2 _03929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05017_ _01504_ _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09825_ _00219_ io_in[4] u_cpu.rf_ram.memory\[43\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09756_ _00150_ io_in[4] u_cpu.rf_ram.memory\[7\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06968_ _02803_ _02827_ _03136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06950__A1 _02766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09802__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08707_ _04266_ _01022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11092__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05919_ _02445_ _02403_ _02446_ _00051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09687_ _04636_ _04832_ _04839_ _01429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06899_ _02891_ _03089_ _03094_ _00385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08298__A4 _03925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08638_ _03922_ _04178_ _04222_ _04225_ _04226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06702__A1 _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08569_ _04164_ _04165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09952__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10600_ _00973_ io_in[4] u_cpu.cpu.decode.op26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07258__A2 _03297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08455__B2 _03901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05269__A1 _01464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10531_ _00904_ io_in[4] u_cpu.rf_ram.memory\[116\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10462_ _00835_ io_in[4] u_cpu.rf_ram.memory\[120\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09000__I _02656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08758__A2 _02598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10393_ _00766_ io_in[4] u_cpu.rf_ram.memory\[36\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05116__S1 _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07430__A2 _03395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09183__A2 _04543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11014_ _01383_ io_in[4] u_cpu.rf_ram.memory\[24\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05744__A2 _02318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06941__A1 _03106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07497__A2 _03425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08446__A1 _03922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07249__A2 _03287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10729_ _01098_ io_in[4] u_cpu.rf_ram.memory\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05680__A1 _01473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05107__S1 _01524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07421__A2 _03385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07940_ _03508_ _03682_ _03689_ _00832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09825__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07871_ _02626_ _02814_ _03651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09610_ u_cpu.rf_ram.memory\[0\]\[4\] _04792_ _04797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08921__A2 _04381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06822_ u_cpu.rf_ram.memory\[68\]\[2\] _03049_ _03052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10802__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05735__A2 _02309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06932__A1 _02827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09541_ _04634_ _04752_ _04758_ _01364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06753_ u_cpu.rf_ram.memory\[74\]\[4\] _03008_ _03013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09975__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05704_ _02259_ _02280_ _02281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09472_ _04622_ _04711_ _04712_ _01341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07488__A2 _03425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06684_ u_cpu.rf_ram.memory\[119\]\[6\] _02967_ _02974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05499__A1 _01465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08423_ _02619_ _02965_ _04040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05635_ u_cpu.rf_ram.memory\[108\]\[7\] u_cpu.rf_ram.memory\[109\]\[7\] u_cpu.rf_ram.memory\[110\]\[7\]
+ u_cpu.rf_ram.memory\[111\]\[7\] _01529_ _01500_ _02213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10952__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06160__A2 _02628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08354_ _02466_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[5\] _03979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05566_ u_cpu.rf_ram.memory\[80\]\[6\] u_cpu.rf_ram.memory\[81\]\[6\] u_cpu.rf_ram.memory\[82\]\[6\]
+ u_cpu.rf_ram.memory\[83\]\[6\] _01544_ _01545_ _02145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_20_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07305_ _03310_ _03325_ _03327_ _00558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08285_ _02465_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[0\] _03913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05497_ _01638_ _02076_ _01534_ _02077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06999__A1 _03110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07236_ u_cpu.rf_ram.memory\[141\]\[7\] _03277_ _03285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07660__A2 _03523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05671__A1 _01465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07167_ _03246_ _03247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06118_ _02265_ u_arbiter.i_wb_cpu_dbus_we _02364_ _02313_ _02604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__07412__A2 _03385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10332__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07098_ u_cpu.rf_ram.memory\[55\]\[1\] _03207_ _03209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05274__I1 u_cpu.rf_ram.memory\[49\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06049_ u_cpu.cpu.ctrl.o_ibus_adr\[23\] u_cpu.cpu.ctrl.o_ibus_adr\[22\] u_cpu.cpu.ctrl.o_ibus_adr\[21\]
+ _02539_ _02548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__04899__I _01485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05974__A2 _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09165__A2 _04533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08912__A2 _04381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09808_ _00202_ io_in[4] u_cpu.rf_ram.memory\[51\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10482__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05726__A2 _02301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09739_ _00133_ io_in[4] u_cpu.rf_ram.memory\[20\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08676__A1 _03697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07479__A2 _03415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08428__A1 _03695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08979__A2 _04425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10514_ _00887_ io_in[4] u_cpu.rf_ram.memory\[122\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05662__A1 _01617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10445_ _00818_ io_in[4] u_cpu.rf_ram.memory\[34\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09848__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07403__A2 _03375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10376_ _00749_ io_in[4] u_cpu.rf_ram.memory\[38\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10825__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09998__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08903__A2 _04371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10975__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06390__A2 _02794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06142__A2 _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10205__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05420_ _01506_ _01999_ _01481_ _02000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05351_ u_cpu.rf_ram.memory\[40\]\[4\] u_cpu.rf_ram.memory\[41\]\[4\] u_cpu.rf_ram.memory\[42\]\[4\]
+ u_cpu.rf_ram.memory\[43\]\[4\] _01551_ _01524_ _01932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__05589__B _01534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08070_ _03701_ _03760_ _03765_ _00886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05282_ _01548_ _01863_ _01579_ _01864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06445__A3 _02622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07642__A2 _03513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10355__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05653__A1 _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07021_ _03114_ _03157_ _03165_ _00436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09395__A2 _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05405__A1 _01966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08972_ _03697_ _04425_ _04428_ _01125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05500__S1 _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09147__A2 _04523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07923_ u_cpu.rf_ram.memory\[34\]\[7\] _03672_ _03680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07854_ u_cpu.cpu.ctrl.i_jump _03611_ _03637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05708__A2 u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06905__A1 _02897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06805_ _02642_ _03039_ _03042_ _00343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07785_ _03502_ _03593_ _03597_ _00768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06381__A2 _02784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04997_ _01565_ _01570_ _01575_ _01580_ _01581_ _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_09524_ u_cpu.cpu.ctrl.i_iscomp _03897_ _04749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06736_ _02891_ _02998_ _03003_ _00313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08658__A1 _03697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09455_ u_cpu.rf_ram.memory\[87\]\[1\] _04701_ _04703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06667_ u_cpu.rf_ram.memory\[40\]\[7\] _02956_ _02964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08406_ _03974_ _04024_ _03938_ _04025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05618_ _01463_ _02195_ _01558_ _02196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11130__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09386_ _04628_ _04661_ _04664_ _01303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07881__A2 _03652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06598_ _02919_ _02921_ _02922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08337_ _03906_ _03917_ _03962_ _03963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05549_ u_cpu.rf_ram.memory\[104\]\[6\] u_cpu.rf_ram.memory\[105\]\[6\] u_cpu.rf_ram.memory\[106\]\[6\]
+ u_cpu.rf_ram.memory\[107\]\[6\] _01555_ _01531_ _02128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_32_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08268_ _03895_ _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07219_ _03114_ _03267_ _03275_ _00524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08199_ u_arbiter.i_wb_cpu_rdt\[14\] _03822_ _03833_ u_arbiter.i_wb_cpu_dbus_dat\[15\]
+ _03853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10848__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__04998__A3 _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09386__A2 _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10230_ _00616_ io_in[4] u_cpu.rf_ram.memory\[137\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07397__A1 _03312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10161_ _00547_ io_in[4] u_cpu.rf_ram.memory\[13\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10092_ _00486_ io_in[4] u_cpu.rf_ram.memory\[53\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10998__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08897__A1 _02642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06372__A2 _02784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10228__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10994_ _01363_ io_in[4] u_cpu.rf_ram.memory\[27\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09310__A2 _04613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07321__A1 _03306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05558__S1 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10378__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07624__A2 _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06017__C _02461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10428_ _00801_ io_in[4] u_cpu.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09377__A2 _04651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10359_ _00019_ io_in[4] u_cpu.rf_ram_if.rdata1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05938__A2 _02456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09129__A2 _04513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05494__S0 _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11003__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04920_ _01504_ _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_78_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04851_ _01438_ u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_54_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06363__A2 _02770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11153__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07570_ _02619_ _02976_ _03474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09301__A2 _04613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06521_ _02742_ _02765_ _02870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_62_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05549__S1 _01531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09240_ _04446_ _04573_ _04579_ _01242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06452_ _02681_ _02829_ _02831_ _00201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05403_ _01977_ _01979_ _01981_ _01983_ _01541_ _01984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_09171_ u_cpu.rf_ram.memory\[104\]\[7\] _04533_ _04541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09065__A1 _04448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06383_ _02689_ _02784_ _02790_ _00173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08122_ _03699_ _03790_ _03794_ _00909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05334_ _01513_ _01914_ _01915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07615__A2 _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08812__A1 u_cpu.cpu.ctrl.o_ibus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08053_ u_cpu.rf_ram.memory\[112\]\[5\] _03750_ _03756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05265_ u_cpu.rf_ram.memory\[44\]\[3\] u_cpu.rf_ram.memory\[45\]\[3\] u_cpu.rf_ram.memory\[46\]\[3\]
+ u_cpu.rf_ram.memory\[47\]\[3\] _01555_ _01531_ _01847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_31_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07004_ _02677_ _02825_ _03156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09368__A2 _04651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05196_ _01512_ _01778_ _01779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07379__A1 _02642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08040__A2 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05485__S0 _01507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08955_ _04403_ _04415_ _03923_ _04416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07906_ _03510_ _03662_ _03670_ _00817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08879__A1 _02642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08886_ u_cpu.rf_ram.memory\[3\]\[6\] _04361_ _04368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_96_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09540__A2 _04752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07837_ u_cpu.rf_ram.memory\[90\]\[1\] _03626_ _03628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06354__A2 _02770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07551__A1 _03322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07768_ u_cpu.rf_ram.memory\[37\]\[4\] _03583_ _03588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04904__A3 _01486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09507_ _01458_ _02302_ _04736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06719_ u_cpu.rf_ram.memory\[139\]\[5\] _02988_ _02994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10520__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07699_ _03506_ _03543_ _03549_ _00730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07303__A1 _03306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08500__B1 _03959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09438_ _04626_ _04691_ _04693_ _01326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07854__A2 _03611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09369_ u_cpu.rf_ram.memory\[10\]\[3\] _04651_ _04655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10670__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06290__A1 _02632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09359__A2 _04641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11026__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10213_ _00599_ io_in[4] u_cpu.rf_ram.memory\[138\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08031__A2 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06042__A1 _02402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05476__S0 _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10144_ _00530_ io_in[4] u_cpu.rf_ram.memory\[141\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10050__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10075_ _00469_ io_in[4] u_cpu.rf_ram.memory\[55\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09531__A2 _04752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08334__A3 _03948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_62_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10977_ _01346_ io_in[4] u_cpu.rf_ram.memory\[88\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08098__A2 _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07845__A2 _03626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09047__A1 u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09598__A2 _04782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05050_ _01622_ _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05084__A2 _01667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08022__A2 _03730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07781__A1 _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08740_ u_arbiter.i_wb_cpu_dbus_adr\[27\] u_arbiter.i_wb_cpu_dbus_adr\[28\] _02335_
+ _04283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05952_ u_cpu.cpu.ctrl.o_ibus_adr\[3\] _02470_ _02471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_85_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05219__S0 _01522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04903_ _01489_ _01490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08671_ u_cpu.rf_ram.memory\[31\]\[0\] _04247_ _04248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10543__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05883_ _02427_ _00032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07533__A1 _03322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06336__A2 _02756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07622_ _03504_ _03496_ _03505_ _00697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07553_ _03464_ _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09286__A1 _04438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08089__A2 _03770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08418__B _03958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06504_ _02860_ _02861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10693__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07836__A2 _03626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07484_ u_cpu.rf_ram.memory\[135\]\[1\] _03425_ _03427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09223_ u_cpu.rf_ram.memory\[105\]\[6\] _04563_ _04570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05847__A1 _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06435_ _02685_ _02816_ _02820_ _00195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09038__A1 _04444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09589__A2 _04782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09154_ _04450_ _04523_ _04531_ _01204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06366_ _02609_ _02673_ _02779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__11049__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08105_ u_cpu.rf_ram.memory\[116\]\[4\] _03780_ _03785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05317_ _01879_ _01898_ _01471_ _01899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09085_ u_arbiter.i_wb_cpu_rdt\[24\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[8\]
+ _04485_ _04494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08261__A2 _03885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06297_ u_cpu.rf_ram.memory\[1\]\[4\] _02733_ _02738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06272__A1 _02683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05075__A2 _01658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08036_ _02657_ _03740_ _03746_ _00871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05248_ _01506_ _01829_ _01519_ _01830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09909__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08013__A2 _03730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10073__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05179_ _01755_ _01757_ _01759_ _01761_ _01560_ _01762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_131_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06024__A1 _02463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09987_ _00381_ io_in[4] u_cpu.rf_ram.memory\[64\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06575__A2 _02900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08938_ _02728_ _04390_ _04400_ _04401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_130_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08869_ _03705_ _04351_ _04358_ _01092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10900_ _01269_ io_in[4] u_cpu.rf_ram.memory\[69\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10831_ _01200_ io_in[4] u_cpu.rf_ram.memory\[103\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__04889__A2 u_cpu.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08328__B _03954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10762_ _01131_ io_in[4] u_cpu.rf_ram.memory\[94\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07827__A2 _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09003__I _02661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05838__A1 _02388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10693_ _01063_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08788__B1 _04311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08252__A2 _03885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10416__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05066__A2 _01649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06263__A1 _01563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08004__A2 _03720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05907__S _02431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10566__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06566__A2 _02731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07763__A1 _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10127_ _00004_ io_in[4] u_cpu.rf_ram.rdata\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10058_ _00452_ io_in[4] u_cpu.rf_ram.memory\[58\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07515__A1 _03322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06318__A2 _02745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09268__A1 _04438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05541__A3 _02119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07818__A2 _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08491__A2 _04093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06220_ _02661_ _02691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06151_ _02611_ u_cpu.rf_ram_if.wdata0_r\[1\] _02634_ _02635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09440__A1 _04628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08243__A2 _03874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10096__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06254__A1 _02685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05102_ _01492_ _01657_ _01666_ _01685_ _01686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_117_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06082_ _02402_ u_scanchain_local.module_data_in\[66\] _02478_ u_arbiter.i_wb_cpu_dbus_adr\[29\]
+ _02575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_99_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10909__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05033_ u_cpu.rf_ram.memory\[84\]\[0\] u_cpu.rf_ram.memory\[85\]\[0\] u_cpu.rf_ram.memory\[86\]\[0\]
+ u_cpu.rf_ram.memory\[87\]\[0\] _01507_ _01605_ _01618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09910_ _00304_ io_in[4] u_cpu.rf_ram.memory\[139\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09841_ _00235_ io_in[4] u_cpu.rf_ram.memory\[47\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08420__C _03965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09772_ _00166_ io_in[4] u_cpu.rf_ram.memory\[78\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_101_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06984_ u_cpu.rf_ram.memory\[61\]\[7\] _03137_ _03145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08723_ _04274_ _01030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05935_ u_arbiter.i_wb_cpu_ibus_adr\[0\] _02456_ _02457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06309__A2 _02745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08654_ _03691_ _04237_ _04238_ _00997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05866_ u_arbiter.i_wb_cpu_rdt\[4\] u_arbiter.i_wb_cpu_dbus_dat\[1\] _02418_ _02419_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_54_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07605_ _02667_ _03485_ _03493_ _00692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08585_ _04000_ _03946_ _03908_ _04177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05797_ _02272_ u_cpu.rf_ram_if.rdata1\[1\] _02370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_35_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07536_ u_cpu.rf_ram.memory\[132\]\[0\] _03455_ _03456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07809__A2 _02259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07467_ _03310_ _03415_ _03417_ _00630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10439__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09206_ _04448_ _04553_ _04560_ _01227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06418_ _02687_ _02805_ _02810_ _00188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07398_ u_cpu.rf_ram.memory\[138\]\[3\] _03375_ _03379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09137_ _02743_ _04349_ _04522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06349_ _02769_ _02770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09731__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08234__A2 _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06245__A1 _02619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09068_ _02910_ _04485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10589__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06796__A2 _03028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08019_ u_cpu.rf_ram.memory\[8\]\[6\] _03730_ _03737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_78_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11030_ _01399_ io_in[4] u_cpu.rf_ram.memory\[98\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09881__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07745__A1 _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05220__A2 _01802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09498__A1 _02305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09498__B2 u_cpu.cpu.state.genblk1.misalign_trap_sync_r vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06720__A2 _02988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10814_ _01183_ io_in[4] u_cpu.rf_ram.memory\[101\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10745_ _01114_ io_in[4] u_cpu.rf_ram.memory\[93\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05287__A2 _01864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10676_ _01048_ io_in[4] u_cpu.rf_ram.memory\[30\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09422__A1 _04628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08225__A2 _03808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06236__A1 _02685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07984__A1 _03705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06787__A2 _03028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06539__A2 _02872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11159_ io_oeb[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_67_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05211__A2 _01793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05720_ _02263_ u_cpu.cpu.genblk3.csr.mcause31 _02292_ _02296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_36_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08161__A1 _02416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05651_ _01464_ _02228_ _02229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06711__A2 _02988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08370_ _03956_ _03992_ _03993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05582_ u_cpu.rf_ram.memory\[128\]\[6\] u_cpu.rf_ram.memory\[129\]\[6\] u_cpu.rf_ram.memory\[130\]\[6\]
+ u_cpu.rf_ram.memory\[131\]\[6\] _01641_ _01635_ _02161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_108_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07321_ _03306_ _03335_ _03336_ _00565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09754__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09661__A1 _04628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06475__A1 _02685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05278__A2 _01831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07252_ u_cpu.rf_ram.memory\[140\]\[6\] _03287_ _03294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06203_ u_cpu.rf_ram.memory\[21\]\[0\] _02679_ _02680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10731__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08216__A2 _03808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07183_ _02667_ _03247_ _03255_ _00508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06227__A1 _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06134_ _02614_ _02618_ _02619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06778__A2 _03018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06065_ u_cpu.cpu.ctrl.o_ibus_adr\[25\] _02561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10881__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05016_ _01597_ _01599_ _01600_ _01601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_132_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07727__A1 _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09824_ _00218_ io_in[4] u_cpu.rf_ram.memory\[43\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10111__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09755_ _00149_ io_in[4] u_cpu.rf_ram.memory\[7\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06967_ _03114_ _03127_ _03135_ _00412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06950__A2 _02827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08706_ u_arbiter.i_wb_cpu_dbus_adr\[10\] u_arbiter.i_wb_cpu_dbus_adr\[11\] _04257_
+ _04266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05918_ u_arbiter.i_wb_cpu_rdt\[29\] _02403_ _02446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09686_ u_cpu.rf_ram.memory\[23\]\[6\] _04832_ _04839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06898_ u_cpu.rf_ram.memory\[64\]\[4\] _03089_ _03094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08152__A1 _03802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08637_ _03955_ _04224_ _04225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05849_ _02406_ _00048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_54_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06702__A2 _02978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10261__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06177__I _02656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08568_ _02259_ _04163_ _02911_ _04164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07519_ _03306_ _03445_ _03446_ _00653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08499_ _03955_ _04101_ _04102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10530_ _00903_ io_in[4] u_cpu.rf_ram.memory\[116\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05269__A2 _01850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06466__A1 _02782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10461_ _00834_ io_in[4] u_cpu.rf_ram.memory\[120\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09404__A1 _04628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08207__A2 _03835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10392_ _00765_ io_in[4] u_cpu.rf_ram.memory\[36\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06769__A2 _03018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05977__B1 _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08341__B _03966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05684__C _01445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11013_ _01382_ io_in[4] u_cpu.rf_ram.memory\[25\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08391__A1 _03936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07194__A2 _03257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08391__B2 _03899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08930__A3 _03948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06941__A2 _03117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04952__A1 _01528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10604__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08143__A1 u_arbiter.i_wb_cpu_dbus_dat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09777__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05920__S _02431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10754__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09643__A1 _04628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10728_ _01097_ io_in[4] u_cpu.rf_ram.memory\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10659_ _01032_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10134__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07709__A1 _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07870_ _02395_ _03602_ _03650_ _00801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08382__A1 _02285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06821_ _02885_ _03049_ _03051_ _00350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05196__A1 _01512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06932__A2 _02870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09540_ u_cpu.rf_ram.memory\[27\]\[5\] _04752_ _04758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05586__I3 u_cpu.rf_ram.memory\[139\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10284__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06752_ _02889_ _03008_ _03012_ _00320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05703_ _02262_ _02278_ _02279_ _02280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09471_ u_cpu.rf_ram.memory\[88\]\[0\] _04711_ _04712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06683_ _02893_ _02967_ _02973_ _00290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_92_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08685__A2 _04247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08422_ _02290_ _03956_ _04039_ _00964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05634_ _01548_ _02211_ _01518_ _02212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05115__B _01600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05499__A2 _02078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06696__A1 _02887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08353_ _03970_ _03971_ _03976_ _03977_ _03978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_51_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05565_ _01597_ _02143_ _01600_ _02144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08437__A2 _04041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04954__B _01482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07304_ u_cpu.rf_ram.memory\[73\]\[1\] _03325_ _03327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08284_ _03904_ _03911_ _03912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05496_ u_cpu.rf_ram.memory\[140\]\[5\] u_cpu.rf_ram.memory\[141\]\[5\] u_cpu.rf_ram.memory\[142\]\[5\]
+ u_cpu.rf_ram.memory\[143\]\[5\] _01634_ _01635_ _02076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_137_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06999__A2 _03147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07235_ _03112_ _03277_ _03284_ _00531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05671__A2 _02248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07166_ _02731_ _02838_ _03246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_117_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06117_ u_cpu.cpu.immdec.imm11_7\[1\] u_cpu.cpu.immdec.imm11_7\[2\] u_cpu.cpu.immdec.imm11_7\[3\]
+ u_cpu.cpu.immdec.imm11_7\[0\] _02603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_07097_ _03098_ _03207_ _03208_ _00469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06048_ u_cpu.cpu.ctrl.o_ibus_adr\[23\] _02546_ _02547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10627__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07176__A2 _03247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08373__A1 _02466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09807_ _00201_ io_in[4] u_cpu.rf_ram.memory\[51\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05187__A1 _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07999_ u_cpu.rf_ram.memory\[121\]\[5\] _03720_ _03726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09738_ _00132_ io_in[4] u_cpu.rf_ram.memory\[20\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07291__I _02656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10777__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09669_ _04636_ _04822_ _04829_ _01421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08676__A2 _04247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06687__A1 _02897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09625__A1 _04628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08428__A2 _04041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04864__B u_cpu.cpu.genblk3.csr.o_new_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10007__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06439__A1 _02689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07100__A2 _03207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10513_ _00886_ io_in[4] u_cpu.rf_ram.memory\[122\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05662__A2 _02239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10444_ _00817_ io_in[4] u_cpu.rf_ram.memory\[35\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10157__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10375_ _00748_ io_in[4] u_cpu.rf_ram.memory\[123\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08600__A2 _04052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08364__A1 _03940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05915__S _02431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05178__A1 _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08116__A1 _03691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08667__A2 _04237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06678__A1 u_cpu.rf_ram.memory\[119\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05350__A1 _01548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06545__I _02636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05350_ _01548_ _01930_ _01518_ _01931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_81_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09092__A2 _04485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05281_ u_cpu.rf_ram.memory\[96\]\[3\] u_cpu.rf_ram.memory\[97\]\[3\] u_cpu.rf_ram.memory\[98\]\[3\]
+ u_cpu.rf_ram.memory\[99\]\[3\] _01567_ _01568_ _01863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__05102__A1 _01492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07020_ u_cpu.rf_ram.memory\[19\]\[7\] _03157_ _03165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11082__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06602__A1 u_cpu.cpu.state.genblk1.misalign_trap_sync_r vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08971_ u_cpu.rf_ram.memory\[97\]\[2\] _04425_ _04428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09942__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07922_ _03508_ _03672_ _03679_ _00824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08355__A1 _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07158__A2 _03237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07853_ _02395_ _03602_ _03635_ _03636_ _00797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__05169__A1 _01513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06905__A2 _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06804_ u_cpu.rf_ram.memory\[6\]\[2\] _03039_ _03042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07784_ u_cpu.rf_ram.memory\[36\]\[3\] _03593_ _03597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04996_ _01485_ _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06735_ u_cpu.rf_ram.memory\[77\]\[4\] _02998_ _03003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09523_ _04747_ _04748_ _01356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08658__A2 _04237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09454_ _04622_ _04701_ _04702_ _01333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06669__A1 _02728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06666_ _02895_ _02956_ _02963_ _00283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07330__A2 _03335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05617_ u_cpu.rf_ram.memory\[44\]\[7\] u_cpu.rf_ram.memory\[45\]\[7\] u_cpu.rf_ram.memory\[46\]\[7\]
+ u_cpu.rf_ram.memory\[47\]\[7\] _01555_ _01531_ _02195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08405_ _03947_ _03972_ _04024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_24_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09385_ u_cpu.rf_ram.memory\[85\]\[2\] _04661_ _04664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05341__A1 _01528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06597_ u_arbiter.i_wb_cpu_dbus_dat\[6\] _02920_ _02921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09607__A1 _02683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08336_ _03906_ _03947_ _03962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05548_ _01512_ _02126_ _02127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07094__A1 _02743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08267_ u_arbiter.i_wb_cpu_ack _02461_ _03894_ _03895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_20_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05479_ _01602_ _02058_ _02059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08830__A2 _04327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07218_ u_cpu.rf_ram.memory\[142\]\[7\] _03267_ _03275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06841__A1 _02887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08198_ u_arbiter.i_wb_cpu_dbus_dat\[14\] _03835_ _03852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07149_ _03236_ _03237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07397__A2 _03375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10160_ _00546_ io_in[4] u_cpu.rf_ram.memory\[13\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10091_ _00485_ io_in[4] u_cpu.rf_ram.memory\[53\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08346__A1 _03922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08897__A2 _04371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04907__A1 _01487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09006__I _02666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10993_ _01362_ io_in[4] u_cpu.rf_ram.memory\[27\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05580__A1 _01492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08649__A2 u_cpu.cpu.genblk3.csr.mstatus_mie vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07321__A2 _03335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05332__A1 _01506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09815__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07085__A1 _03106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05191__S0 _01551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09965__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10427_ _00800_ io_in[4] u_cpu.cpu.bufreg2.i_cnt_done vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08585__A1 _04000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05709__I _01441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07388__A2 _03365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10358_ _00018_ io_in[4] u_cpu.rf_ram_if.rdata1\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10942__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05494__S1 _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10289_ _00675_ io_in[4] u_cpu.rf_ram.memory\[131\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08337__A1 _03906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08888__A2 _04361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04850_ _01437_ _01438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06899__A1 _02891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07560__A2 _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06520_ _02693_ _02861_ _02869_ _00231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_18_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07312__A2 _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06451_ u_cpu.rf_ram.memory\[51\]\[1\] _02829_ _02831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10322__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05323__A1 _01465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05402_ _01617_ _01982_ _01481_ _01983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_21_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09170_ _04448_ _04533_ _04540_ _01211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06382_ u_cpu.rf_ram.memory\[42\]\[5\] _02784_ _02790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09065__A2 _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08121_ u_cpu.rf_ram.memory\[33\]\[3\] _03790_ _03794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05333_ u_cpu.rf_ram.memory\[20\]\[4\] u_cpu.rf_ram.memory\[21\]\[4\] u_cpu.rf_ram.memory\[22\]\[4\]
+ u_cpu.rf_ram.memory\[23\]\[4\] _01497_ _01501_ _01914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07076__A1 _02827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08812__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10472__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08052_ _03701_ _03750_ _03755_ _00878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06823__A1 _02887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05264_ _01505_ _01845_ _01846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05182__S0 _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07003_ _03114_ _03147_ _03155_ _00428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05195_ u_cpu.rf_ram.memory\[108\]\[2\] u_cpu.rf_ram.memory\[109\]\[2\] u_cpu.rf_ram.memory\[110\]\[2\]
+ u_cpu.rf_ram.memory\[111\]\[2\] _01529_ _01524_ _01778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_116_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07379__A2 _03365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06051__A2 _02397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08954_ _03903_ _03918_ _04031_ _04415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05485__S1 _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07905_ u_cpu.rf_ram.memory\[35\]\[7\] _03662_ _03670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08879__A2 _04361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08885_ _02657_ _04361_ _04367_ _01099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_96_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07836_ _03494_ _03626_ _03627_ _00789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07551__A2 _03455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04979_ u_cpu.rf_ram.memory\[60\]\[0\] u_cpu.rf_ram.memory\[61\]\[0\] u_cpu.rf_ram.memory\[62\]\[0\]
+ u_cpu.rf_ram.memory\[63\]\[0\] _01562_ _01563_ _01564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_71_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07767_ _03502_ _03583_ _03587_ _00760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04904__A4 _01490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09506_ _04732_ _04723_ _04735_ _02302_ _01352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_53_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06718_ _02891_ _02988_ _02993_ _00305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09838__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07698_ u_cpu.rf_ram.memory\[125\]\[5\] _03543_ _03549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07303__A2 _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08500__B2 _04099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09437_ u_cpu.rf_ram.memory\[111\]\[1\] _04691_ _04693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05314__A1 _01512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06649_ _02897_ _02945_ _02953_ _00276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10815__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09368_ _02642_ _04651_ _04654_ _01295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_40_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09056__A2 _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07067__A1 _03106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06118__C _02313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09988__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08319_ u_arbiter.i_wb_cpu_rdt\[15\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\]
+ _02465_ _03947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09299_ _02675_ _02768_ _04612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08614__B _03924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05173__S0 _01495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10965__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06290__A2 _02733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08567__A1 _01444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10212_ _00598_ io_in[4] u_cpu.rf_ram.memory\[138\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10143_ _00529_ io_in[4] u_cpu.rf_ram.memory\[141\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05476__S1 _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07790__A2 _03593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10074_ _00468_ io_in[4] u_cpu.rf_ram.memory\[56\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07542__A2 _03455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10345__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05553__A1 _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09295__A2 _04603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10976_ _01345_ io_in[4] u_cpu.rf_ram.memory\[88\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05305__A1 _01617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10495__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05213__B _01600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07058__A1 _02827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06805__A1 _02642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05164__S0 _01530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06281__A2 _02719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08558__A1 _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11120__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07781__A2 _03593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05951_ _02467_ u_cpu.cpu.ctrl.o_ibus_adr\[2\] _02470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04902_ _01487_ _01488_ _01489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_78_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08670_ _04246_ _04247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05219__S1 _01622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05882_ u_arbiter.i_wb_cpu_rdt\[12\] u_arbiter.i_wb_cpu_dbus_dat\[9\] _02418_ _02427_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07533__A2 _03445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07621_ u_cpu.rf_ram.memory\[22\]\[4\] _03496_ _03505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05544__A1 _01512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07552_ _02825_ _02976_ _03464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10838__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09286__A2 _04603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06503_ _02754_ _02827_ _02860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07483_ _03306_ _03425_ _03426_ _00637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08494__B1 _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09222_ _04446_ _04563_ _04569_ _01234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06434_ u_cpu.rf_ram.memory\[44\]\[3\] _02816_ _02820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05847__A2 _02355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09038__A2 _04463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09153_ u_cpu.rf_ram.memory\[103\]\[7\] _04523_ _04531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07049__A1 _03106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06365_ _02693_ _02770_ _02778_ _00167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08246__B1 _03874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10988__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08104_ _03699_ _03780_ _03784_ _00901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05316_ _01492_ _01888_ _01897_ _01898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_09084_ _04493_ _01172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05155__S0 _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06296_ _02647_ _02733_ _02737_ _00139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08035_ u_cpu.rf_ram.memory\[11\]\[5\] _03740_ _03746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06272__A2 _02719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05247_ u_cpu.rf_ram.memory\[16\]\[3\] u_cpu.rf_ram.memory\[17\]\[3\] u_cpu.rf_ram.memory\[18\]\[3\]
+ u_cpu.rf_ram.memory\[19\]\[3\] _01508_ _01509_ _01829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_135_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10218__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05178_ _01554_ _01760_ _01558_ _01761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09986_ _00380_ io_in[4] u_cpu.rf_ram.memory\[65\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07772__A2 _03583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10368__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08937_ u_cpu.cpu.immdec.imm11_7\[1\] _04390_ _04400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08868_ u_cpu.rf_ram.memory\[109\]\[6\] _04351_ _04358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07524__A2 _03445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07819_ u_cpu.rf_ram.memory\[91\]\[1\] _03616_ _03618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05535__A1 _01548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08799_ _04319_ _01061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_10830_ _01199_ io_in[4] u_cpu.rf_ram.memory\[103\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09277__A2 _04593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10761_ _01130_ io_in[4] u_cpu.rf_ram.memory\[97\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08485__B1 _03909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05838__A2 _02397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09029__A2 _04463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10692_ _01062_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08237__B1 _03829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05146__S0 _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11143__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09201__A2 _04553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08960__A1 _04024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10126_ _00003_ io_in[4] u_cpu.rf_ram.rdata\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07763__A2 _03583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05774__A1 _01441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10057_ _00451_ io_in[4] u_cpu.rf_ram.memory\[58\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07515__A2 _03435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05526__A1 _01504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09268__A2 _04593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08476__B1 _04075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10959_ _01328_ io_in[4] u_cpu.rf_ram.memory\[111\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08779__A1 _03707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06150_ _02606_ u_cpu.rf_ram_if.wdata1_r\[1\] _02634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_129_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05137__S0 _01529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09440__A2 _04691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05101_ _01490_ _01675_ _01684_ _01685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__06254__A2 _02707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06081_ u_cpu.cpu.ctrl.o_ibus_adr\[29\] _02571_ _02574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07451__A1 _03312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05032_ _01463_ _01617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10510__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09840_ _00234_ io_in[4] u_cpu.rf_ram.memory\[47\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07754__A2 _03573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09771_ _00165_ io_in[4] u_cpu.rf_ram.memory\[78\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05765__A1 _02336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06983_ _03112_ _03137_ _03144_ _00419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08722_ u_arbiter.i_wb_cpu_dbus_adr\[18\] u_arbiter.i_wb_cpu_dbus_adr\[19\] _02335_
+ _04274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05934_ _02455_ _02456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10660__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07506__A2 _03435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08653_ u_cpu.rf_ram.memory\[32\]\[0\] _04237_ _04238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05865_ _02388_ _02418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05517__A1 _01528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07604_ u_cpu.rf_ram.memory\[12\]\[7\] _03485_ _03493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_42_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09259__A2 _04583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08584_ _03910_ _03985_ _04150_ _04176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05796_ _02273_ u_cpu.rf_ram.rdata\[1\] _02369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06190__A1 u_cpu.rf_ram.memory\[82\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11016__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07535_ _03454_ _03455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07466_ u_cpu.rf_ram.memory\[136\]\[1\] _03415_ _03417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05376__S0 _01496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09205_ u_cpu.rf_ram.memory\[79\]\[6\] _04553_ _04560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06417_ u_cpu.rf_ram.memory\[45\]\[4\] _02805_ _02810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06493__A2 _02851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07397_ _03312_ _03375_ _03378_ _00599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10040__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09136_ _04450_ _04513_ _04521_ _01196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06348_ _02766_ _02768_ _02769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05128__S0 _01507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09431__A2 _04681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06245__A2 _02677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09067_ _04450_ _04476_ _04484_ _01164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06279_ u_cpu.rf_ram.memory\[20\]\[6\] _02719_ _02726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07993__A2 _03720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08018_ _02657_ _03730_ _03736_ _00863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_78_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10190__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07294__I _02661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08942__A1 _03924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07745__A2 _03573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09969_ _00363_ io_in[4] u_cpu.rf_ram.memory\[67\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05300__S0 _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09498__A2 _02400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05508__A1 _01506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06181__A1 _02611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10813_ _01182_ io_in[4] u_cpu.rf_ram.memory\[101\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10744_ _01113_ io_in[4] u_cpu.rf_ram.memory\[93\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05367__S0 _01551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09670__A2 _04822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07681__A1 _03506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10675_ _01047_ io_in[4] u_cpu.rf_ram.memory\[30\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09422__A2 _04681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10533__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07433__A1 _03312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06236__A2 _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07984__A2 _03710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09186__A1 _04446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10683__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07736__A2 _03563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08933__A1 _03910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11158_ io_oeb[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_96_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05747__A1 _02263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10109_ _00503_ io_in[4] u_cpu.rf_ram.memory\[9\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11089_ _00037_ io_in[0] u_arbiter.i_wb_cpu_ack vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11039__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08161__A2 _03822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05650_ u_cpu.rf_ram.memory\[92\]\[7\] u_cpu.rf_ram.memory\[93\]\[7\] u_cpu.rf_ram.memory\[94\]\[7\]
+ u_cpu.rf_ram.memory\[95\]\[7\] _01562_ _01563_ _02228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_63_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06548__I _02641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06172__A1 u_cpu.rf_ram.memory\[82\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05581_ _02140_ _02159_ _01471_ _02160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10063__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09110__A1 _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07320_ u_cpu.rf_ram.memory\[71\]\[0\] _03335_ _03336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05358__S0 _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09661__A2 _04822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07251_ _03110_ _03287_ _03293_ _00538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06475__A2 _02840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05278__A3 _01840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06202_ _02678_ _02679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06283__I u_cpu.cpu.immdec.imm11_7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07182_ u_cpu.rf_ram.memory\[9\]\[7\] _03247_ _03255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09413__A2 _04671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06133_ _01500_ _02617_ _02618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05120__C _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06227__A2 _02695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07975__A2 _03710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06064_ u_cpu.cpu.ctrl.o_ibus_adr\[26\] _02560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05986__A1 _02463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05015_ _01480_ _01600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07727__A2 _03563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09823_ _00217_ io_in[4] u_cpu.rf_ram.memory\[43\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09754_ _00148_ io_in[4] u_cpu.rf_ram.memory\[7\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06966_ u_cpu.rf_ram.memory\[62\]\[7\] _03127_ _03135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08705_ _04265_ _01021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05917_ u_arbiter.i_wb_cpu_dbus_dat\[26\] _02445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09685_ _04634_ _04832_ _04838_ _01428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06897_ _02889_ _03089_ _03093_ _00384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08636_ _02467_ u_arbiter.i_wb_cpu_rdt\[19\] _03912_ _04223_ _04224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__10406__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05848_ u_arbiter.i_wb_cpu_ack _02389_ _02405_ _02406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06163__A1 _02611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05597__S0 _01530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08567_ _01444_ _02328_ _02269_ _02318_ _04163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_54_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05779_ _02285_ u_cpu.cpu.mem_bytecnt\[1\] _02291_ _02282_ _02354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09101__A1 _02675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07518_ u_cpu.rf_ram.memory\[133\]\[0\] _03445_ _03446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08498_ _02265_ _04100_ _02392_ _04101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_70_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05349__S0 _01495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09652__A2 _04812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10556__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07663__A1 _03506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08606__C _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06466__A2 _02838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07449_ _03310_ _03405_ _03407_ _00622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_7_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10460_ _00833_ io_in[4] u_cpu.rf_ram.memory\[117\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09404__A2 _04671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09119_ _03037_ _04349_ _04512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06218__A2 _02679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07415__A1 _03312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10391_ _00764_ io_in[4] u_cpu.rf_ram.memory\[37\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05977__A1 _02403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09168__A1 _04446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08915__A1 _03697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07718__A2 _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11012_ _01381_ io_in[4] u_cpu.rf_ram.memory\[25\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05981__B _02456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08930__A4 _03962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04952__A2 _01536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10086__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08143__A2 _02915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05588__S0 _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09643__A2 _04812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08446__A3 _04000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10727_ _01096_ io_in[4] u_cpu.rf_ram.memory\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06457__A2 _02829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08851__B1 _04329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10658_ _01031_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06209__A2 _02679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10589_ _00962_ io_in[4] u_cpu.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07709__A2 _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08382__A2 _03956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06820_ u_cpu.rf_ram.memory\[68\]\[1\] _03049_ _03051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10429__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05196__A2 _01778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06393__A1 _02681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06751_ u_cpu.rf_ram.memory\[74\]\[3\] _03008_ _03012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09721__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05702_ u_cpu.cpu.alu.i_rs1 u_cpu.cpu.alu.add_cy_r _02279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09470_ _04710_ _04711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06682_ u_cpu.rf_ram.memory\[119\]\[5\] _02967_ _02973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08694__S _04257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10579__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08421_ _03965_ _04030_ _04038_ _03955_ _04039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05633_ u_cpu.rf_ram.memory\[96\]\[7\] u_cpu.rf_ram.memory\[97\]\[7\] u_cpu.rf_ram.memory\[98\]\[7\]
+ u_cpu.rf_ram.memory\[99\]\[7\] _01567_ _01568_ _02211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_52_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06696__A2 _02978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05564_ u_cpu.rf_ram.memory\[88\]\[6\] u_cpu.rf_ram.memory\[89\]\[6\] u_cpu.rf_ram.memory\[90\]\[6\]
+ u_cpu.rf_ram.memory\[91\]\[6\] _01598_ _01556_ _02143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08352_ _03963_ _03977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09634__A2 _04802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09871__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07303_ _03306_ _03325_ _03326_ _00557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07645__A1 _03506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08842__B1 _04329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08283_ _03909_ _03910_ _03911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05495_ _01465_ _02074_ _02075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07234_ u_cpu.rf_ram.memory\[141\]\[6\] _03277_ _03284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07165_ _03114_ _03237_ _03245_ _00500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06116_ _01460_ _01456_ _02392_ u_cpu.cpu.o_wen1 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08070__A1 _03701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07096_ u_cpu.rf_ram.memory\[55\]\[0\] _03207_ _03208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05959__A1 _02464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06047_ u_cpu.cpu.ctrl.o_ibus_adr\[22\] u_cpu.cpu.ctrl.o_ibus_adr\[21\] _02539_ _02546_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_59_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06620__A2 _02935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09806_ _00200_ io_in[4] u_cpu.rf_ram.memory\[51\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05187__A2 _01769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07998_ _03701_ _03720_ _03725_ _00854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09737_ _00131_ io_in[4] u_cpu.rf_ram.memory\[20\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06949_ _03114_ _03117_ _03125_ _00404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08125__A2 _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09668_ u_cpu.rf_ram.memory\[89\]\[6\] _04822_ _04829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08619_ u_cpu.cpu.immdec.imm19_12_20\[7\] _03955_ _04209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07884__A1 _03506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06687__A2 _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09599_ _04638_ _04782_ _04790_ _01390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_54_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09625__A2 _04802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04864__C u_cpu.cpu.state.genblk1.misalign_trap_sync_r vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06439__A2 _02816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07636__A1 u_cpu.rf_ram.memory\[128\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10512_ _00885_ io_in[4] u_cpu.rf_ram.memory\[122\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05041__B _01519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05111__A2 _01690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10443_ _00816_ io_in[4] u_cpu.rf_ram.memory\[35\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04870__A1 _01444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07939__A2 _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10374_ _00747_ io_in[4] u_cpu.rf_ram.memory\[123\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08600__A3 _04111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09744__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09561__A1 _04636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08364__A2 _03941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06375__A1 _02681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10721__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08116__A2 _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06127__A1 u_cpu.cpu.immdec.imm11_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09894__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06678__A2 _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10871__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05730__I _01445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09616__A2 _04792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05350__A2 _01930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07627__A1 u_cpu.rf_ram.memory\[22\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08824__B1 _04329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05280_ _01571_ _01861_ _01862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05102__A2 _01657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10101__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06850__A2 _03059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08052__A1 _03701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08970_ _03695_ _04425_ _04427_ _01124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10251__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07921_ u_cpu.rf_ram.memory\[34\]\[6\] _03672_ _03679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08355__A2 u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07852_ u_cpu.cpu.state.genblk1.misalign_trap_sync_r _03611_ _03636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06803_ _02637_ _03039_ _03041_ _00342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_84_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07783_ _03500_ _03593_ _03596_ _00767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_49_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_04995_ _01505_ _01578_ _01579_ _01580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08107__A2 _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09304__A1 _04438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09522_ u_cpu.cpu.genblk3.csr.mstatus_mie _04720_ _04745_ _04748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06734_ _02889_ _02998_ _03002_ _00312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06118__A1 _02265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09453_ u_cpu.rf_ram.memory\[87\]\[0\] _04701_ _04702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06665_ u_cpu.rf_ram.memory\[40\]\[6\] _02956_ _02963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04965__B _01518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08404_ _03901_ _04022_ _04023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05616_ _01505_ _02193_ _02194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09384_ _04626_ _04661_ _04663_ _01302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06596_ _02263_ _02598_ _02314_ _02920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05341__A2 _01921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09607__A2 _04792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07618__A1 u_cpu.rf_ram.memory\[22\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08335_ _03914_ _03906_ _03961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05547_ u_cpu.rf_ram.memory\[108\]\[6\] u_cpu.rf_ram.memory\[109\]\[6\] u_cpu.rf_ram.memory\[110\]\[6\]
+ u_cpu.rf_ram.memory\[111\]\[6\] _01529_ _01500_ _02126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08815__B1 _04311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08266_ _02909_ u_arbiter.i_wb_cpu_ibus_adr\[1\] _03894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08291__A1 _03906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07094__A2 _02827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05478_ u_cpu.rf_ram.memory\[80\]\[5\] u_cpu.rf_ram.memory\[81\]\[5\] u_cpu.rf_ram.memory\[82\]\[5\]
+ u_cpu.rf_ram.memory\[83\]\[5\] _01544_ _01545_ _02058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07217_ _03112_ _03267_ _03274_ _00523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06841__A2 _03059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08197_ _03850_ _03851_ _00927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07148_ _02717_ _02827_ _03236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09767__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07079_ _03098_ _03197_ _03198_ _00461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10090_ _00484_ io_in[4] u_cpu.rf_ram.memory\[54\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10744__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09543__A1 _04636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08346__A2 _03923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06357__A1 _02685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04907__A2 _01488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10894__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10992_ _01361_ io_in[4] u_cpu.rf_ram.memory\[27\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08649__A3 u_cpu.cpu.genblk3.csr.i_mtip vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07857__A1 _02277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05332__A2 _01912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10124__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07609__A1 u_cpu.rf_ram.memory\[22\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08806__B1 _04311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07085__A2 _03197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08282__A1 _03901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06832__A2 _03049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10274__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05191__S1 _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05891__I0 u_arbiter.i_wb_cpu_rdt\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08034__A1 _02652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10426_ _00799_ io_in[4] u_cpu.cpu.ctrl.i_jump vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06045__B1 _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10357_ _00017_ io_in[4] u_cpu.rf_ram_if.rdata1\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06596__A1 _02263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10288_ _00674_ io_in[4] u_cpu.rf_ram.memory\[131\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08337__A2 _03917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06348__A1 _02766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06899__A2 _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07848__A1 _03508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06450_ _02669_ _02829_ _02830_ _00200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06520__A1 _02693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05401_ u_cpu.rf_ram.memory\[76\]\[4\] u_cpu.rf_ram.memory\[77\]\[4\] u_cpu.rf_ram.memory\[78\]\[4\]
+ u_cpu.rf_ram.memory\[79\]\[4\] _01529_ _01500_ _01982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_61_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06381_ _02687_ _02784_ _02789_ _00172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05332_ _01506_ _01912_ _01481_ _01913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08120_ _03697_ _03790_ _03793_ _00908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10617__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07076__A2 _02954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08051_ u_cpu.rf_ram.memory\[112\]\[4\] _03750_ _03755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05263_ u_cpu.rf_ram.memory\[40\]\[3\] u_cpu.rf_ram.memory\[41\]\[3\] u_cpu.rf_ram.memory\[42\]\[3\]
+ u_cpu.rf_ram.memory\[43\]\[3\] _01551_ _01524_ _01845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06823__A2 _03049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05182__S1 _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05882__I0 u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07002_ u_cpu.rf_ram.memory\[60\]\[7\] _03147_ _03155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05194_ _01548_ _01776_ _01579_ _01777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09073__I0 u_arbiter.i_wb_cpu_rdt\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10767__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08576__A2 _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06587__A1 u_cpu.cpu.state.genblk1.misalign_trap_sync_r vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08953_ u_cpu.cpu.immdec.imm11_7\[3\] _04390_ _03897_ _04414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08328__A2 _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09525__A1 _03966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07904_ _03508_ _03662_ _03669_ _00816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08884_ u_cpu.rf_ram.memory\[3\]\[5\] _04361_ _04367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06339__A1 _02689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07835_ u_cpu.rf_ram.memory\[90\]\[0\] _03626_ _03627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07000__A2 _03147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05011__A1 _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07766_ u_cpu.rf_ram.memory\[37\]\[3\] _03583_ _03587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04978_ _01499_ _01563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10147__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09505_ _02325_ _04725_ _04723_ _04735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_25_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06717_ u_cpu.rf_ram.memory\[139\]\[4\] _02988_ _02993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07697_ _03504_ _03543_ _03548_ _00729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08500__A2 _03956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09436_ _04622_ _04691_ _04692_ _01325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06648_ u_cpu.rf_ram.memory\[17\]\[7\] _02945_ _02953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05314__A2 _01895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09367_ u_cpu.rf_ram.memory\[10\]\[2\] _04651_ _04654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06579_ _02657_ _02900_ _02906_ _00253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10297__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08318_ _03942_ _03944_ _03945_ _03899_ _03946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__07067__A2 _03187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09298_ _04450_ _04603_ _04611_ _01268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08249_ _03884_ _03885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06814__A2 _03039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07297__I _02666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05173__S1 _01499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08016__A1 _02652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10211_ _00597_ io_in[4] u_cpu.rf_ram.memory\[138\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10142_ _00528_ io_in[4] u_cpu.rf_ram.memory\[141\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09516__A1 _02293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10073_ _00467_ io_in[4] u_cpu.rf_ram.memory\[56\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06750__A1 _02887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11072__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10975_ _01344_ io_in[4] u_cpu.rf_ram.memory\[88\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05305__A2 _01886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06502__A1 _02693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09932__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09047__A3 _02461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08255__A1 _03697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07058__A2 _02838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06805__A2 _03039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05164__S1 _01532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10409_ _00782_ io_in[4] u_cpu.rf_ram.memory\[91\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06569__A1 _02632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07230__A2 _03277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05950_ _02469_ _00060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_61_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04901_ u_cpu.cpu.immdec.imm24_20\[3\] _01469_ _01488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05881_ _02426_ _00031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07620_ _02651_ _03504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_94_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07551_ _03322_ _03455_ _03463_ _00668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06502_ _02693_ _02851_ _02859_ _00223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08494__A1 _03935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07482_ u_cpu.rf_ram.memory\[135\]\[0\] _03425_ _03426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08494__B2 _03961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09221_ u_cpu.rf_ram.memory\[105\]\[5\] _04563_ _04569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06433_ _02683_ _02816_ _02819_ _00194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09152_ _04448_ _04523_ _04530_ _01203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07049__A2 _03177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08246__A1 u_arbiter.i_wb_cpu_rdt\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06364_ u_cpu.rf_ram.memory\[78\]\[7\] _02770_ _02778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08246__B2 _02277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08103_ u_cpu.rf_ram.memory\[116\]\[3\] _03780_ _03784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05315_ _01890_ _01892_ _01894_ _01896_ _01541_ _01897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_09083_ u_arbiter.i_wb_cpu_rdt\[23\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[7\]
+ _04485_ _04493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06295_ u_cpu.rf_ram.memory\[1\]\[3\] _02733_ _02737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05155__S1 _01509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08034_ _02652_ _03740_ _03745_ _00870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05246_ _01513_ _01827_ _01828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08549__A2 _02585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05177_ u_cpu.rf_ram.memory\[44\]\[2\] u_cpu.rf_ram.memory\[45\]\[2\] u_cpu.rf_ram.memory\[46\]\[2\]
+ u_cpu.rf_ram.memory\[47\]\[2\] _01555_ _01531_ _01760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_118_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09985_ _00379_ io_in[4] u_cpu.rf_ram.memory\[65\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08936_ _03956_ _04398_ _04399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09805__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11095__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08867_ _03703_ _04351_ _04357_ _01091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07818_ _03494_ _03616_ _03617_ _00781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_17_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06732__A1 _02887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08798_ u_cpu.cpu.ctrl.o_ibus_adr\[7\] _04309_ _04311_ u_cpu.cpu.ctrl.o_ibus_adr\[8\]
+ _04319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_77_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07749_ _03502_ _03573_ _03577_ _00752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09955__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05314__B _01481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10760_ _01129_ io_in[4] u_cpu.rf_ram.memory\[97\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08485__A1 _03922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08485__B2 _04088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05299__A1 _01464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09419_ u_cpu.rf_ram.memory\[86\]\[1\] _04681_ _04683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10932__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10691_ _01061_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08237__A1 u_arbiter.i_wb_cpu_rdt\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08237__B2 u_arbiter.i_wb_cpu_dbus_dat\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08788__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05146__S1 _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07460__A2 _03405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05471__A1 _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07212__A2 _03267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10312__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10125_ _00002_ io_in[4] u_cpu.rf_ram.rdata\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05774__A2 _02309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06971__A1 _03098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10056_ _00450_ io_in[4] u_cpu.rf_ram.memory\[58\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05208__C _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10462__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06723__A1 u_cpu.rf_ram.memory\[139\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05526__A2 _02104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08476__A1 _03941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10958_ _01327_ io_in[4] u_cpu.rf_ram.memory\[111\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08476__B2 _03947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10889_ _01258_ io_in[4] u_cpu.rf_ram.memory\[83\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08779__A2 _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05137__S1 _01500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05100_ _01677_ _01679_ _01681_ _01683_ _01581_ _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_06080_ _02570_ _02572_ _02573_ _00088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07451__A2 _03405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05462__A1 _01566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05031_ _01602_ _01615_ _01616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09828__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09770_ _00164_ io_in[4] u_cpu.rf_ram.memory\[78\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06982_ u_cpu.rf_ram.memory\[61\]\[6\] _03137_ _03144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10805__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08721_ _04273_ _01029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05933_ _02401_ _02397_ _02455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_113_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09978__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08652_ _04236_ _04237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_94_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05864_ _02416_ _02389_ _02417_ _00092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05517__A2 _02095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06714__A1 _02887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04957__C _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07603_ _02662_ _03485_ _03492_ _00691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_81_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08583_ _04149_ _04174_ _04175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10955__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05795_ _02368_ u_cpu.cpu.o_wdata0 vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_35_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06190__A2 _02628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05134__B _01519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07534_ _02717_ _02976_ _03454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07465_ _03306_ _03415_ _03416_ _00629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05376__S1 _01594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09204_ _04446_ _04553_ _04559_ _01226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06416_ _02685_ _02805_ _02809_ _00187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08219__A1 u_arbiter.i_wb_cpu_dbus_dat\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07690__A2 _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07396_ u_cpu.rf_ram.memory\[138\]\[2\] _03375_ _03378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09135_ u_cpu.rf_ram.memory\[102\]\[7\] _04513_ _04521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06347_ _02767_ _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05128__S1 _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09066_ u_cpu.rf_ram.memory\[28\]\[7\] _04476_ _04484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06278_ _02689_ _02719_ _02725_ _00133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07442__A2 _03395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10335__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05453__A1 _01490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08017_ u_cpu.rf_ram.memory\[8\]\[5\] _03730_ _03736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05229_ _01792_ _01811_ _01471_ _01812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_78_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09195__A2 _04553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05205__A1 _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09968_ _00362_ io_in[4] u_cpu.rf_ram.memory\[67\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10485__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05300__S1 _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06953__A1 _03098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08919_ _03701_ _04381_ _04386_ _01114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09899_ _00293_ io_in[4] u_cpu.rf_ram.memory\[129\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05508__A2 _02086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06181__A2 u_cpu.rf_ram_if.wdata0_r\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10812_ _01181_ io_in[4] u_cpu.rf_ram.memory\[101\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08458__A1 _04009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10743_ _01112_ io_in[4] u_cpu.rf_ram.memory\[93\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07130__A1 _02675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05367__S1 _01524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11110__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07681__A2 _03533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10674_ _01046_ io_in[4] u_cpu.rf_ram.memory\[30\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05692__A1 _01444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08630__A1 u_cpu.cpu.immdec.imm19_12_20\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07433__A2 _03395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05995__A2 _02397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10828__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09186__A2 _04543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07197__A1 _02657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11157_ _00091_ io_in[0] u_scanchain_local.module_data_in\[69\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05747__A2 _02320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10108_ _00502_ io_in[4] u_cpu.rf_ram.memory\[9\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11088_ _00026_ io_in[0] u_cpu.cpu.genblk3.csr.i_mtip vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10978__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10039_ _00433_ io_in[4] u_cpu.rf_ram.memory\[19\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06172__A2 _02628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10208__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08449__A1 _04000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05580_ _01492_ _02149_ _02158_ _02159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_17_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09110__A2 _04503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07121__A1 _03106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05358__S1 _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07250_ u_cpu.rf_ram.memory\[140\]\[5\] _03287_ _03293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07672__A2 _03533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10358__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06201_ _02675_ _02677_ _02678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05683__A1 _01441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07181_ _02662_ _03247_ _03254_ _00507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06132_ _02616_ _02617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_129_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08621__A1 _03959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07424__A2 _03385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06063_ _02463_ _02558_ _02559_ _00085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09177__A2 _04543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05014_ u_cpu.rf_ram.memory\[120\]\[0\] u_cpu.rf_ram.memory\[121\]\[0\] u_cpu.rf_ram.memory\[122\]\[0\]
+ u_cpu.rf_ram.memory\[123\]\[0\] _01598_ _01556_ _01599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_28_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09822_ _00216_ io_in[4] u_cpu.rf_ram.memory\[43\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08924__A2 _04381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05129__B _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06935__A1 _03098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05294__S0 _01576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09753_ _00147_ io_in[4] u_cpu.rf_ram.memory\[7\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06965_ _03112_ _03127_ _03134_ _00411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08704_ u_arbiter.i_wb_cpu_dbus_adr\[9\] u_arbiter.i_wb_cpu_dbus_adr\[10\] _04257_
+ _04265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05916_ _02444_ _00050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09684_ u_cpu.rf_ram.memory\[23\]\[5\] _04832_ _04838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08688__A1 _02392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06896_ u_cpu.rf_ram.memory\[64\]\[3\] _03089_ _03093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08635_ _02467_ _02416_ _04223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05847_ _02306_ _02355_ _02388_ _02405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05597__S1 _01532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11133__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08566_ _04160_ _04161_ _04162_ _03897_ _00985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05778_ u_cpu.cpu.mem_if.signbit _02353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_70_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09101__A2 _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07517_ _03444_ _03445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_126_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08497_ _01444_ _02305_ u_arbiter.i_wb_cpu_dbus_we _04100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__07112__A1 _02827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05349__S1 _01499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07448_ u_cpu.rf_ram.memory\[49\]\[1\] _03405_ _03407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07663__A2 _03523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07379_ _02642_ _03365_ _03368_ _00591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_136_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09118_ _04450_ _04503_ _04511_ _01188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08612__A1 _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10390_ _00763_ io_in[4] u_cpu.rf_ram.memory\[37\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07415__A2 _03385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09049_ _02395_ _04474_ _01156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_2_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09168__A2 _04533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07179__A1 _02657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11011_ _01380_ io_in[4] u_cpu.rf_ram.memory\[25\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08915__A2 _04381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05285__S0 _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06154__A2 _02628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07351__A1 _03320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05588__S1 _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10500__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07103__A1 _03106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08446__A4 _03998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10726_ _01095_ io_in[4] u_cpu.rf_ram.memory\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07654__A2 _03523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08851__B2 _04347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10657_ _01030_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10650__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08603__A1 _04031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07406__A2 _03375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10588_ _00961_ io_in[4] u_cpu.cpu.csr_d_sel vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09159__A2 _04533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11006__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06052__C _02388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08906__A2 _04371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07943__I _02631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06393__A2 _02794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11156__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10030__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06750_ _02887_ _03008_ _03011_ _00319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_77_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05028__S0 _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05701_ _02261_ _02277_ _02278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_37_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06681_ _02891_ _02967_ _02972_ _00289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06145__A2 _02611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08390__I0 u_arbiter.i_wb_cpu_rdt\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08420_ _04031_ _04032_ _04037_ _03965_ _04038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_36_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05632_ _01512_ _02209_ _02210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07893__A2 _03662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10180__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08351_ _03926_ _03928_ _03972_ _03975_ _03976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05563_ _01464_ _02141_ _02142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07302_ u_cpu.rf_ram.memory\[73\]\[0\] _03325_ _03326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08282_ _03901_ _03903_ _03910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05494_ u_cpu.rf_ram.memory\[136\]\[5\] u_cpu.rf_ram.memory\[137\]\[5\] u_cpu.rf_ram.memory\[138\]\[5\]
+ u_cpu.rf_ram.memory\[139\]\[5\] _01634_ _01635_ _02074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07645__A2 _03513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05200__S0 _01496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07233_ _03110_ _03277_ _03283_ _00530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07164_ u_cpu.rf_ram.memory\[52\]\[7\] _03237_ _03245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06115_ _02600_ _02602_ _02599_ _00023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_133_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08070__A2 _03760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07095_ _03206_ _03207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06046_ _02463_ _02544_ _02545_ _00082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09570__A2 _04772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09805_ _00199_ io_in[4] u_cpu.rf_ram.memory\[44\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07997_ u_cpu.rf_ram.memory\[121\]\[4\] _03720_ _03725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07581__A1 _03316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06384__A2 _02784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09736_ _00130_ io_in[4] u_cpu.rf_ram.memory\[20\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06948_ u_cpu.rf_ram.memory\[63\]\[7\] _03117_ _03125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10523__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09667_ _04634_ _04822_ _04828_ _01420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06879_ _02889_ _03079_ _03083_ _00376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05306__C _01486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07333__A1 _03320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08618_ _04206_ _04207_ _04159_ _04208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07884__A2 _03652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09598_ u_cpu.rf_ram.memory\[24\]\[7\] _04782_ _04790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08617__C _04031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08549_ u_cpu.cpu.immdec.imm7 _02585_ _04106_ _04146_ _04147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_42_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10673__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07636__A2 _03513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05647__A1 _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10511_ _00884_ io_in[4] u_cpu.rf_ram.memory\[122\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09389__A2 _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10442_ _00815_ io_in[4] u_cpu.rf_ram.memory\[35\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11029__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04870__A2 _01445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10373_ _00746_ io_in[4] u_cpu.rf_ram.memory\[123\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08061__A2 _03760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10053__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09561__A2 _04762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06375__A2 _02784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09313__A2 _04613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06127__A2 _02611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07875__A2 _03652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05430__S0 _01523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07627__A2 _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05638__A1 _01566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10709_ _01079_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05102__A3 _01666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08052__A2 _03750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06063__A1 _02463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05810__A1 _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07920_ _03506_ _03672_ _03678_ _00823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09552__A2 _04762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07851_ _01444_ _02305_ _02391_ _03635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__10546__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07563__A1 _03316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06802_ u_cpu.rf_ram.memory\[6\]\[1\] _03039_ _03041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07782_ u_cpu.rf_ram.memory\[36\]\[2\] _03593_ _03596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04994_ _01518_ _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09521_ _01477_ _02301_ _04746_ _04747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06733_ u_cpu.rf_ram.memory\[77\]\[3\] _02998_ _03002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09304__A2 _04613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06118__A2 u_arbiter.i_wb_cpu_dbus_we vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07315__A1 _03320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09452_ _04700_ _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10696__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06664_ _02893_ _02956_ _02962_ _00282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08403_ _04000_ _03930_ _04022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05421__S0 _01497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05615_ u_cpu.rf_ram.memory\[40\]\[7\] u_cpu.rf_ram.memory\[41\]\[7\] u_cpu.rf_ram.memory\[42\]\[7\]
+ u_cpu.rf_ram.memory\[43\]\[7\] _01551_ _01524_ _02193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09383_ u_cpu.rf_ram.memory\[85\]\[1\] _04661_ _04663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06595_ _02915_ _02918_ _02919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08334_ _03936_ _03938_ _03948_ _03960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_05546_ _01548_ _02124_ _01579_ _02125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07618__A2 _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08265_ _03707_ _03885_ _03893_ _00953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05477_ _01597_ _02056_ _01600_ _02057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08291__A2 _03908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07216_ u_cpu.rf_ram.memory\[142\]\[6\] _03267_ _03274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08196_ u_arbiter.i_wb_cpu_rdt\[13\] _03822_ _03833_ u_arbiter.i_wb_cpu_dbus_dat\[14\]
+ _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_134_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07147_ _03114_ _03227_ _03235_ _00492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09240__A1 _04446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08043__A2 _03750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10076__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07078_ u_cpu.rf_ram.memory\[56\]\[0\] _03197_ _03198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05801__A1 _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06029_ _02461_ _02530_ _02531_ _02532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_133_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09543__A2 _04752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06357__A2 _02770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05317__B _01471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09719_ _00113_ io_in[4] u_cpu.rf_ram.memory\[81\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10991_ _01360_ io_in[4] u_cpu.rf_ram.memory\[27\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05580__A3 _02158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08628__B _03965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05412__S0 _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09059__A1 _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07609__A2 _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08282__A2 _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10419__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10425_ _00798_ io_in[4] u_cpu.cpu.mem_if.signbit vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09711__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08034__A2 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06045__A1 _02402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08585__A3 _03908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10356_ _00016_ io_in[4] u_cpu.rf_ram_if.rdata1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10569__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06596__A2 _02598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07793__A1 _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10287_ _00673_ io_in[4] u_cpu.rf_ram.memory\[131\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09861__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09534__A2 _04752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04910__I _01494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06348__A2 _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07545__A1 _03316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09298__A1 _04450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07848__A2 _03626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06058__B _02397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06520__A2 _02861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05400_ _01621_ _01980_ _01981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06380_ u_cpu.rf_ram.memory\[42\]\[4\] _02784_ _02789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05331_ u_cpu.rf_ram.memory\[24\]\[4\] u_cpu.rf_ram.memory\[25\]\[4\] u_cpu.rf_ram.memory\[26\]\[4\]
+ u_cpu.rf_ram.memory\[27\]\[4\] _01508_ _01509_ _01912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_119_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10099__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08050_ _03699_ _03750_ _03754_ _00877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06284__A1 u_cpu.cpu.immdec.imm11_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05262_ _01548_ _01843_ _01518_ _01844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_31_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07001_ _03112_ _03147_ _03154_ _00427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05193_ u_cpu.rf_ram.memory\[96\]\[2\] u_cpu.rf_ram.memory\[97\]\[2\] u_cpu.rf_ram.memory\[98\]\[2\]
+ u_cpu.rf_ram.memory\[99\]\[2\] _01567_ _01568_ _01776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09222__A1 _04446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08025__A2 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06036__A1 _02463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08952_ u_cpu.cpu.immdec.imm11_7\[4\] _02392_ _02604_ _04413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_102_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07903_ u_cpu.rf_ram.memory\[35\]\[6\] _03662_ _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08883_ _02652_ _04361_ _04366_ _01098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_111_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06339__A2 _02756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07834_ _03625_ _03626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05011__A2 _01595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05642__S0 _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07765_ _03500_ _03583_ _03586_ _00759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_04977_ _01495_ _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_65_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09504_ _04734_ _01351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06716_ _02889_ _02988_ _02992_ _00304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07839__A2 _03626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07696_ u_cpu.rf_ram.memory\[125\]\[4\] _03543_ _03548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09435_ u_cpu.rf_ram.memory\[111\]\[0\] _04691_ _04692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06647_ _02895_ _02945_ _02952_ _00275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06511__A2 _02861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09366_ _02637_ _04651_ _04653_ _01294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_36_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06578_ u_cpu.rf_ram.memory\[4\]\[5\] _02900_ _02906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08317_ u_arbiter.i_wb_cpu_rdt\[4\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[4\]
+ _02466_ _03945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05529_ u_cpu.rf_ram.memory\[44\]\[6\] u_cpu.rf_ram.memory\[45\]\[6\] u_cpu.rf_ram.memory\[46\]\[6\]
+ u_cpu.rf_ram.memory\[47\]\[6\] _01555_ _01531_ _02108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09297_ u_cpu.rf_ram.memory\[108\]\[7\] _04603_ _04611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08264__A2 _03885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09734__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08248_ _02695_ _02965_ _03884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05600__B _01519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10711__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08016__A2 _03730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08179_ _03838_ _03839_ _00921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10210_ _00596_ io_in[4] u_cpu.rf_ram.memory\[14\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09884__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06578__A2 _02900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07775__A1 _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10141_ _00527_ io_in[4] u_cpu.rf_ram.memory\[141\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10861__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09516__A2 _03605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10072_ _00466_ io_in[4] u_cpu.rf_ram.memory\[56\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07527__A1 _03316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05633__S0 _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08358__B _03982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06750__A2 _03008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10974_ _01343_ io_in[4] u_cpu.rf_ram.memory\[88\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08488__C1 _04088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06502__A2 _02851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10241__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08255__A2 _03885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10391__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09204__A1 _04446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08007__A2 _03730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10408_ _00781_ io_in[4] u_cpu.rf_ram.memory\[91\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08313__S _02465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06569__A2 _02900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08540__C _03998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10339_ _00725_ io_in[4] u_cpu.rf_ram.memory\[125\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04900_ u_cpu.cpu.immdec.imm19_12_20\[7\] _01438_ _01487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05880_ u_arbiter.i_wb_cpu_rdt\[11\] u_arbiter.i_wb_cpu_dbus_dat\[8\] _02418_ _02426_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_66_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07951__I _02641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05624__S0 _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06741__A2 _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07550_ u_cpu.rf_ram.memory\[132\]\[7\] _03455_ _03463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06501_ u_cpu.rf_ram.memory\[43\]\[7\] _02851_ _02859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07481_ _03424_ _03425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08494__A2 _03914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09757__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09220_ _04444_ _04563_ _04568_ _01233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06432_ u_cpu.rf_ram.memory\[44\]\[2\] _02816_ _02819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09151_ u_cpu.rf_ram.memory\[103\]\[6\] _04523_ _04530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06363_ _02691_ _02770_ _02777_ _00166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10734__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08246__A2 _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08102_ _03697_ _03780_ _03783_ _00900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05314_ _01512_ _01895_ _01481_ _01896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05420__B _01481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09082_ _04492_ _01171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06294_ _02642_ _02733_ _02736_ _00138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08033_ u_cpu.rf_ram.memory\[11\]\[4\] _03740_ _03745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05245_ u_cpu.rf_ram.memory\[20\]\[3\] u_cpu.rf_ram.memory\[21\]\[3\] u_cpu.rf_ram.memory\[22\]\[3\]
+ u_cpu.rf_ram.memory\[23\]\[3\] _01497_ _01501_ _01827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_116_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10884__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05176_ _01505_ _01758_ _01759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07757__A1 _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09984_ _00378_ io_in[4] u_cpu.rf_ram.memory\[65\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08935_ _04393_ _04396_ _04397_ _03910_ _04398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10114__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07509__A1 _03316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06980__A2 _03137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08866_ u_cpu.rf_ram.memory\[109\]\[5\] _04351_ _04357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05615__S0 _01551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07817_ u_cpu.rf_ram.memory\[91\]\[0\] _03616_ _03617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08797_ _04318_ _01060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_72_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06732__A2 _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10264__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07748_ u_cpu.rf_ram.memory\[38\]\[3\] _03573_ _03577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07679_ _03504_ _03533_ _03538_ _00721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08485__A2 _03908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05299__A2 _01880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06496__A1 _02687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09418_ _04622_ _04681_ _04682_ _01317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_16_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10690_ _01060_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08625__C _03915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08237__A2 _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09349_ u_cpu.rf_ram.memory\[59\]\[2\] _04641_ _04644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06248__A1 _02669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07996__A1 _03699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06015__A4 u_cpu.cpu.ctrl.o_ibus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06420__A1 _02689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10124_ _00001_ io_in[4] u_cpu.rf_ram.rdata\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06971__A2 _03137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10055_ _00449_ io_in[4] u_cpu.rf_ram.memory\[58\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10607__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05606__S0 _01497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06723__A2 _02988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07920__A1 _03506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10757__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10957_ _01326_ io_in[4] u_cpu.rf_ram.memory\[111\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08476__A2 _04051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10888_ _01257_ io_in[4] u_cpu.rf_ram.memory\[83\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08228__A2 _03833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07987__A1 _02838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05030_ u_cpu.rf_ram.memory\[80\]\[0\] u_cpu.rf_ram.memory\[81\]\[0\] u_cpu.rf_ram.memory\[82\]\[0\]
+ u_cpu.rf_ram.memory\[83\]\[0\] _01496_ _01594_ _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10137__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07739__A1 _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08400__A2 _03956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06981_ _03110_ _03137_ _03143_ _00418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06962__A2 _03127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08720_ u_arbiter.i_wb_cpu_dbus_adr\[17\] u_arbiter.i_wb_cpu_dbus_adr\[18\] _04257_
+ _04273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05932_ _02403_ u_scanchain_local.module_data_in\[37\] _02454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10287__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08164__A1 _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08651_ _02754_ _02782_ _04236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05863_ u_arbiter.i_wb_cpu_dbus_dat\[0\] _02389_ _02417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06714__A2 _02988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07602_ u_cpu.rf_ram.memory\[12\]\[6\] _03485_ _03492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08582_ _03980_ _03976_ _04173_ _04052_ _04174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05794_ _01460_ _02343_ _02352_ _02367_ _02368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_07533_ _03322_ _03445_ _03453_ _00660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07464_ u_cpu.rf_ram.memory\[136\]\[0\] _03415_ _03416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09203_ u_cpu.rf_ram.memory\[79\]\[5\] _04553_ _04559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06415_ u_cpu.rf_ram.memory\[45\]\[3\] _02805_ _02809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08219__A2 _03808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07395_ _03310_ _03375_ _03377_ _00598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09134_ _04448_ _04513_ _04520_ _01195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06346_ _02728_ _02608_ _02623_ _02729_ _02767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_136_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07978__A1 _03699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09065_ _04448_ _04476_ _04483_ _01163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06277_ u_cpu.rf_ram.memory\[20\]\[5\] _02719_ _02725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08016_ _02652_ _03730_ _03735_ _00862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05228_ _01492_ _01801_ _01810_ _01811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__05453__A2 _02023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11062__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05159_ u_cpu.rf_ram.memory\[16\]\[2\] u_cpu.rf_ram.memory\[17\]\[2\] u_cpu.rf_ram.memory\[18\]\[2\]
+ u_cpu.rf_ram.memory\[19\]\[2\] _01508_ _01509_ _01742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__05205__A2 _01787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09967_ _00361_ io_in[4] u_cpu.rf_ram.memory\[67\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06953__A2 _03127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09922__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08918_ u_cpu.rf_ram.memory\[93\]\[4\] _04381_ _04386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09898_ _00292_ io_in[4] u_cpu.rf_ram.memory\[119\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08849_ _02276_ _02334_ _01451_ _04346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_57_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06705__A2 _02978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07902__A1 _03506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05325__B _01534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10811_ _01180_ io_in[4] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08458__A2 _04050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08636__B _03912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06469__A1 _02669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10742_ _01111_ io_in[4] u_cpu.rf_ram.memory\[93\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07130__A2 _02827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05141__A1 _01705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10673_ _01045_ io_in[4] u_cpu.cpu.bufreg.lsb\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05692__A2 _01445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07969__A1 _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08371__B _03993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08630__A2 _03955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06641__A1 _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08394__A1 _03901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07197__A2 _03257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11156_ _00090_ io_in[0] u_scanchain_local.module_data_in\[68\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06944__A2 _03117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10107_ _00501_ io_in[4] u_cpu.rf_ram.memory\[9\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11087_ u_scanchain_local.module_data_in\[69\] io_in[0] u_scanchain_local.data_out
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_49_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08146__A1 u_arbiter.i_wb_cpu_dbus_dat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10038_ _00432_ io_in[4] u_cpu.rf_ram.memory\[19\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08449__A2 _03929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07121__A2 _03217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05132__A1 _01621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06200_ _02676_ _02677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05683__A2 u_cpu.cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07180_ u_cpu.rf_ram.memory\[9\]\[6\] _03247_ _03254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11085__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06131_ _01494_ _02615_ _02616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_118_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08621__A2 _04202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06632__A1 _02677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06062_ _02402_ u_scanchain_local.module_data_in\[62\] _02478_ u_arbiter.i_wb_cpu_dbus_adr\[25\]
+ _02559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_144_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05013_ _01495_ _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09945__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08385__A1 _04000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07188__A2 _03257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08385__B2 _03945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09821_ _00215_ io_in[4] u_cpu.rf_ram.memory\[41\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06935__A2 _03117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10922__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05294__S1 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09752_ _00146_ io_in[4] u_cpu.rf_ram.memory\[7\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_101_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06964_ u_cpu.rf_ram.memory\[62\]\[6\] _03127_ _03134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08137__A1 u_arbiter.i_wb_cpu_dbus_dat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08703_ _04264_ _01020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_104_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05915_ u_arbiter.i_wb_cpu_rdt\[28\] u_arbiter.i_wb_cpu_dbus_dat\[25\] _02431_ _02444_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_27_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09683_ _04632_ _04832_ _04837_ _01427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06895_ _02887_ _03089_ _03092_ _00383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05846_ _02400_ _02398_ _02404_ _00037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08634_ _04013_ _04221_ _03969_ _04222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05145__B _01482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07360__A2 _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08565_ u_cpu.cpu.immdec.imm7 _02259_ _04162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05777_ _02313_ _02305_ _02265_ _02351_ _02352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_39_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07516_ _02675_ _02976_ _03444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08496_ u_arbiter.i_wb_cpu_rdt\[25\] u_arbiter.i_wb_cpu_rdt\[9\] _02467_ _04099_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_120_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07112__A2 _03037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10302__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05123__A1 _01464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07447_ _03306_ _03405_ _03406_ _00621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08860__A2 _04351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07378_ u_cpu.rf_ram.memory\[14\]\[2\] _03365_ _03368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_109_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09117_ u_cpu.rf_ram.memory\[101\]\[7\] _04503_ _04511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06329_ _02669_ _02756_ _02757_ _00152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08612__A2 _02411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10452__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06623__A1 _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09048_ _02467_ _04473_ _04474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_124_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11010_ _01379_ io_in[4] u_cpu.rf_ram.memory\[25\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07179__A2 _03247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05285__S1 _01531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08128__A1 _03705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08679__A2 _04247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05055__B _01534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07351__A2 _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09818__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08300__A1 _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07103__A2 _03207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10725_ _01094_ io_in[4] u_cpu.rf_ram.memory\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05502__C _01466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10656_ _01029_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09968__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08603__A2 _03961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10587_ _00960_ io_in[4] u_cpu.cpu.decode.co_mem_word vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06614__A1 _02677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10945__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11139_ _00072_ io_in[0] u_scanchain_local.module_data_in\[51\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07590__A2 _03485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05700_ _02271_ _02276_ u_arbiter.i_wb_cpu_dbus_we _02277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__05028__S1 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06680_ u_cpu.rf_ram.memory\[119\]\[4\] _02967_ _02972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07342__A2 _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05631_ u_cpu.rf_ram.memory\[100\]\[7\] u_cpu.rf_ram.memory\[101\]\[7\] u_cpu.rf_ram.memory\[102\]\[7\]
+ u_cpu.rf_ram.memory\[103\]\[7\] _01551_ _01524_ _02209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_92_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10325__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08390__I1 u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08350_ _03974_ _03947_ _03975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05562_ u_cpu.rf_ram.memory\[92\]\[6\] u_cpu.rf_ram.memory\[93\]\[6\] u_cpu.rf_ram.memory\[94\]\[6\]
+ u_cpu.rf_ram.memory\[95\]\[6\] _01562_ _01563_ _02141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_51_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07301_ _03324_ _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08281_ _03906_ _03908_ _03909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05493_ _02053_ _02072_ _01471_ _02073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08842__A2 _04327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10475__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07232_ u_cpu.rf_ram.memory\[141\]\[5\] _03277_ _03283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05200__S1 _01594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07163_ _03112_ _03237_ _03244_ _00499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06114_ _02601_ _02362_ _02602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07094_ _02743_ _02827_ _03206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06045_ _02402_ u_scanchain_local.module_data_in\[59\] _02478_ u_arbiter.i_wb_cpu_dbus_adr\[22\]
+ _02545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08358__A1 _02400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09804_ _00198_ io_in[4] u_cpu.rf_ram.memory\[44\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07996_ _03699_ _03720_ _03724_ _00853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11100__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07581__A2 _03475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09735_ _00129_ io_in[4] u_cpu.rf_ram.memory\[20\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06947_ _03112_ _03117_ _03124_ _00403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05592__A1 _01473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09666_ u_cpu.rf_ram.memory\[89\]\[5\] _04822_ _04828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06878_ u_cpu.rf_ram.memory\[65\]\[3\] _03079_ _03083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07333__A2 _03335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08617_ _03924_ _03906_ _03909_ _04202_ _04031_ _04207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05829_ _02388_ _02389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09597_ _04636_ _04782_ _04789_ _01389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10818__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08548_ _04143_ _04144_ _04145_ _02585_ _04146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_70_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07097__A1 _03098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08479_ u_cpu.cpu.immdec.imm24_20\[4\] _03955_ _04084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10510_ _00883_ io_in[4] u_cpu.rf_ram.memory\[122\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10968__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10441_ _00814_ io_in[4] u_cpu.rf_ram.memory\[35\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08597__A1 _03972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05829__I _02388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10372_ _00745_ io_in[4] u_cpu.rf_ram.memory\[123\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06072__A2 _02562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08349__A1 _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07021__A1 _03114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07572__A2 _03475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10348__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05583__A1 _01465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07324__A2 _03335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10498__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05430__S1 _01525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04908__I _01464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09790__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08824__A2 _04327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10708_ _01078_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10639_ _01012_ io_in[4] u_cpu.rf_ram.memory\[31\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__04941__S0 _01523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08588__A1 _03908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07954__I _02646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11123__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09001__A2 _04436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07850_ _03510_ _03626_ _03634_ _00796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07563__A2 _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06801_ _02632_ _03039_ _03040_ _00341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_68_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05574__A1 _01617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04993_ u_cpu.rf_ram.memory\[48\]\[0\] u_cpu.rf_ram.memory\[49\]\[0\] u_cpu.rf_ram.memory\[50\]\[0\]
+ u_cpu.rf_ram.memory\[51\]\[0\] _01576_ _01577_ _01578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07781_ _03498_ _03593_ _03595_ _00766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09520_ _04739_ _01477_ _02303_ _04745_ _04746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_06732_ _02887_ _02998_ _03001_ _00311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07315__A2 _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09451_ _02626_ _02743_ _04700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06663_ u_cpu.rf_ram.memory\[40\]\[5\] _02956_ _02962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08402_ _03944_ _03988_ _04021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05614_ _01504_ _02191_ _01518_ _02192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05421__S1 _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09382_ _04622_ _04661_ _04662_ _01301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06594_ u_arbiter.i_wb_cpu_dbus_dat\[5\] _02917_ _02918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_80_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07079__A1 _03098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05545_ u_cpu.rf_ram.memory\[96\]\[6\] u_cpu.rf_ram.memory\[97\]\[6\] u_cpu.rf_ram.memory\[98\]\[6\]
+ u_cpu.rf_ram.memory\[99\]\[6\] _01567_ _01568_ _02124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08333_ _02911_ _03912_ _03959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08815__A2 _04327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08264_ u_cpu.rf_ram.memory\[113\]\[7\] _03885_ _03893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05629__A2 _02197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05476_ u_cpu.rf_ram.memory\[88\]\[5\] u_cpu.rf_ram.memory\[89\]\[5\] u_cpu.rf_ram.memory\[90\]\[5\]
+ u_cpu.rf_ram.memory\[91\]\[5\] _01598_ _01556_ _02056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_20_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07215_ _03110_ _03267_ _03273_ _00522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08195_ u_arbiter.i_wb_cpu_dbus_dat\[13\] _03835_ _03850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07146_ u_cpu.rf_ram.memory\[53\]\[7\] _03227_ _03235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09240__A2 _04573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07251__A1 _03110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07077_ _03196_ _03197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06028_ u_cpu.cpu.ctrl.o_ibus_adr\[19\] u_cpu.cpu.ctrl.o_ibus_adr\[18\] _02508_ _02520_
+ _02531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_82_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05801__A2 _02371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07003__A1 _03114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08751__A1 _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07554__A2 _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05565__A1 _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07979_ u_cpu.rf_ram.memory\[118\]\[4\] _03710_ _03715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09718_ _00112_ io_in[4] u_cpu.rf_ram.memory\[81\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10990_ _01359_ io_in[4] u_cpu.rf_ram.memory\[27\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10640__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07306__A2 _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09649_ _04634_ _04812_ _04818_ _01412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05317__A1 _01879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05412__S1 _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09059__A2 _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10790__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08806__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06293__A2 _02733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10020__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11146__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10424_ _00797_ io_in[4] u_cpu.cpu.state.genblk1.misalign_trap_sync_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09231__A2 _04573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10355_ _00015_ io_in[4] u_cpu.rf_ram_if.rdata1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08990__A1 _04438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07793__A2 _03593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10286_ _00672_ io_in[4] u_cpu.rf_ram.memory\[131\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10170__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05508__B _01481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07545__A2 _03455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05227__C _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09298__A2 _04603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05308__A1 _01621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05330_ _01493_ _01910_ _01911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06853__I _03068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05261_ u_cpu.rf_ram.memory\[32\]\[3\] u_cpu.rf_ram.memory\[33\]\[3\] u_cpu.rf_ram.memory\[34\]\[3\]
+ u_cpu.rf_ram.memory\[35\]\[3\] _01495_ _01499_ _01843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_30_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06284__A2 _02608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06074__B _02402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07000_ u_cpu.rf_ram.memory\[60\]\[6\] _03147_ _03154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05192_ _01571_ _01774_ _01775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09222__A2 _04563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10513__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07233__A1 _03110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07784__A2 _03593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08951_ _04404_ _04410_ _04412_ _01120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07902_ _03506_ _03662_ _03668_ _00815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08882_ u_cpu.rf_ram.memory\[3\]\[4\] _04361_ _04366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10663__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07536__A2 _03455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07833_ _02626_ _02780_ _03625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05642__S1 _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07764_ u_cpu.rf_ram.memory\[37\]\[2\] _03583_ _03586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09289__A2 _04603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04976_ _01547_ _01550_ _01553_ _01559_ _01560_ _01561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__11019__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04976__C _01560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09503_ _04733_ u_cpu.cpu.genblk3.csr.mcause3_0\[2\] _04723_ _04734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_53_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06715_ u_cpu.rf_ram.memory\[139\]\[3\] _02988_ _02992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07695_ _03502_ _03543_ _03547_ _00728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_92_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09434_ _04690_ _04691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06646_ u_cpu.rf_ram.memory\[17\]\[6\] _02945_ _02952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09365_ u_cpu.rf_ram.memory\[10\]\[1\] _04651_ _04653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06577_ _02652_ _02900_ _02905_ _00252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10043__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08316_ _02465_ _02416_ _03943_ _03944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05528_ _01505_ _02106_ _02107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09296_ _04448_ _04603_ _04610_ _01267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09461__A2 _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05459_ u_cpu.rf_ram.memory\[108\]\[5\] u_cpu.rf_ram.memory\[109\]\[5\] u_cpu.rf_ram.memory\[110\]\[5\]
+ u_cpu.rf_ram.memory\[111\]\[5\] _01529_ _01500_ _02039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06275__A2 _02719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08247_ _02452_ _03835_ _03883_ _00945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_21_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08178_ u_arbiter.i_wb_cpu_rdt\[7\] _03822_ _03833_ u_arbiter.i_wb_cpu_dbus_dat\[8\]
+ _03839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10193__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09213__A2 _04563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08272__I0 u_arbiter.i_wb_cpu_rdt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07129_ _03114_ _03217_ _03225_ _00484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08972__A1 _03697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10140_ _00526_ io_in[4] u_cpu.rf_ram.memory\[141\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07775__A2 _03583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10071_ _00465_ io_in[4] u_cpu.rf_ram.memory\[56\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07527__A2 _03445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08639__B _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05633__S1 _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05842__I _02388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08488__B1 _04070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10973_ _01342_ io_in[4] u_cpu.rf_ram.memory\[88\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08488__C2 _04009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05397__S0 _01507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10536__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09204__A2 _04553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06018__A2 _02397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07215__A1 _03110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10407_ _00780_ io_in[4] u_cpu.cpu.state.o_cnt_r\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10686__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08963__A1 u_cpu.cpu.immdec.imm30_25\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07766__A2 _03583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04921__I _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10338_ _00724_ io_in[4] u_cpu.rf_ram.memory\[126\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05777__A1 _02313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10269_ _00655_ io_in[4] u_cpu.rf_ram.memory\[133\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07518__A2 _03445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08549__B _04106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05624__S1 _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05752__I _02265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09140__A1 _04434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10066__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06500_ _02691_ _02851_ _02858_ _00222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07480_ _02743_ _02976_ _03424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05388__S0 _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06431_ _02681_ _02816_ _02818_ _00193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09150_ _04446_ _04523_ _04529_ _01202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06362_ u_cpu.rf_ram.memory\[78\]\[6\] _02770_ _02777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09443__A2 _04691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05313_ u_cpu.rf_ram.memory\[76\]\[3\] u_cpu.rf_ram.memory\[77\]\[3\] u_cpu.rf_ram.memory\[78\]\[3\]
+ u_cpu.rf_ram.memory\[79\]\[3\] _01529_ _01500_ _01895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08101_ u_cpu.rf_ram.memory\[116\]\[2\] _03780_ _03783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06257__A2 _02707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07454__A1 u_cpu.rf_ram.memory\[49\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09081_ u_arbiter.i_wb_cpu_rdt\[22\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[6\]
+ _04485_ _04492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06293_ u_cpu.rf_ram.memory\[1\]\[2\] _02733_ _02736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05244_ _01506_ _01825_ _01481_ _01826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08032_ _02647_ _03740_ _03744_ _00869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06009__A2 u_cpu.cpu.ctrl.o_ibus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05175_ u_cpu.rf_ram.memory\[40\]\[2\] u_cpu.rf_ram.memory\[41\]\[2\] u_cpu.rf_ram.memory\[42\]\[2\]
+ u_cpu.rf_ram.memory\[43\]\[2\] _01551_ _01524_ _01758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07757__A2 _03573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08954__A1 _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05768__A1 _02305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09983_ _00377_ io_in[4] u_cpu.rf_ram.memory\[65\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08934_ _03944_ _03908_ _03909_ _03932_ _04397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_112_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07509__A2 _03435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08865_ _03701_ _04351_ _04356_ _01090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08459__B _04067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07816_ _03615_ _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10409__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05615__S1 _01524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08796_ u_cpu.cpu.ctrl.o_ibus_adr\[6\] _04309_ _04311_ u_cpu.cpu.ctrl.o_ibus_adr\[7\]
+ _04318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_45_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07747_ _03500_ _03573_ _03576_ _00751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05940__A1 _02396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04959_ _01495_ _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07678_ u_cpu.rf_ram.memory\[126\]\[4\] _03533_ _03538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09682__A2 _04832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09417_ u_cpu.rf_ram.memory\[86\]\[0\] _04681_ _04682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10559__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07693__A1 _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06496__A2 _02851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06629_ _02895_ _02935_ _02942_ _00267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_12_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09348_ _04626_ _04641_ _04643_ _01286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09851__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06248__A2 _02707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09279_ u_cpu.rf_ram.memory\[83\]\[7\] _04593_ _04601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07996__A2 _03720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09198__A1 _04440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07748__A2 _03573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05759__A1 u_cpu.cpu.state.o_cnt_r\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06420__A2 _02805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10123_ _00000_ io_in[4] u_cpu.rf_ram.rdata\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10054_ _00448_ io_in[4] u_cpu.rf_ram.memory\[58\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09370__A1 _02647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10089__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05606__S1 _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06184__A1 u_cpu.rf_ram.memory\[82\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07920__A2 _03672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09122__A1 _04434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10956_ _01325_ io_in[4] u_cpu.rf_ram.memory\[111\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06487__A2 _02851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10887_ _01256_ io_in[4] u_cpu.rf_ram.memory\[83\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05521__B _01482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04916__I _01500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09425__A2 _04681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06239__A2 _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08484__I0 u_arbiter.i_wb_cpu_rdt\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07987__A2 _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07739__A2 _03563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08936__A1 _03956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06411__A2 _02805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06980_ u_cpu.rf_ram.memory\[61\]\[5\] _03137_ _03143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05931_ _02452_ _02403_ _02453_ _00056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09724__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08164__A2 _03802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09361__A1 _02731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08650_ _04233_ _04234_ _04235_ _00996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_93_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05862_ u_arbiter.i_wb_cpu_rdt\[3\] _02416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06175__A1 _02611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07601_ _02657_ _03485_ _03491_ _00690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07911__A2 _03672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08581_ _04000_ _03918_ _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10701__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05793_ _02305_ _02318_ _02341_ _02366_ _02367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_82_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07532_ u_cpu.rf_ram.memory\[133\]\[7\] _03445_ _03453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09874__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09664__A2 _04822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07675__A1 _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07463_ _03414_ _03415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06478__A2 _02840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09202_ _04444_ _04553_ _04558_ _01225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06414_ _02683_ _02805_ _02808_ _00186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10851__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07394_ u_cpu.rf_ram.memory\[138\]\[1\] _03375_ _03377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05781__S0 _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09133_ u_cpu.rf_ram.memory\[102\]\[6\] _04513_ _04520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05150__C _01466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06345_ _02618_ _02765_ _02766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_120_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07978__A2 _03710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06276_ _02687_ _02719_ _02724_ _00132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09064_ u_cpu.rf_ram.memory\[28\]\[6\] _04476_ _04483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05227_ _01803_ _01805_ _01807_ _01809_ _01541_ _01810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_08015_ u_cpu.rf_ram.memory\[8\]\[4\] _03730_ _03735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05453__A3 _02032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08927__A1 _03955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05158_ _01513_ _01740_ _01741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06402__A2 _02794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09966_ _00360_ io_in[4] u_cpu.rf_ram.memory\[67\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05089_ u_cpu.rf_ram.memory\[44\]\[1\] u_cpu.rf_ram.memory\[45\]\[1\] u_cpu.rf_ram.memory\[46\]\[1\]
+ u_cpu.rf_ram.memory\[47\]\[1\] _01555_ _01531_ _01673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10231__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08917_ _03699_ _04381_ _04385_ _01113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09897_ _00291_ io_in[4] u_cpu.rf_ram.memory\[119\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09352__A1 _04630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08155__A2 _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08848_ _02363_ _02341_ u_cpu.cpu.ctrl.i_jump _04345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_57_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07902__A2 _03662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10381__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08779_ _03707_ _04299_ _04307_ _01053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09104__A1 _04434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10810_ _01179_ io_in[4] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10741_ _01110_ io_in[4] u_cpu.rf_ram.memory\[93\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06469__A2 _02840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05341__B _01534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10672_ _01044_ io_in[4] u_cpu.cpu.bufreg.lsb\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09407__A2 _04671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05692__A3 _01442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07969__A2 _03037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06641__A2 _02945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09747__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09591__A1 _04630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11155_ _00089_ io_in[0] u_scanchain_local.module_data_in\[67\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05601__B1 _02176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10106_ _00500_ io_in[4] u_cpu.rf_ram.memory\[52\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11086_ u_cpu.cpu.o_wen1 io_in[4] u_cpu.rf_ram_if.wen1_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10724__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09343__A1 _02827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10037_ _00431_ io_in[4] u_cpu.rf_ram.memory\[19\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06157__A1 _02611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09897__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10874__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08319__S _02465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09646__A2 _04812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07657__A1 _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10939_ _01308_ io_in[4] u_cpu.rf_ram.memory\[85\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05132__A2 _01715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10104__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06880__A2 _03079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07957__I _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04891__A1 _01438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06130_ u_cpu.rf_ram_if.rcnt\[0\] u_cpu.rf_ram_if.rcnt\[1\] u_cpu.rf_ram_if.rcnt\[2\]
+ _02615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08082__A1 _03695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06061_ u_cpu.cpu.ctrl.o_ibus_adr\[25\] _02554_ _02558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06632__A2 _02695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10254__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05012_ _01504_ _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09582__A1 _02677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08385__A2 _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09820_ _00214_ io_in[4] u_cpu.rf_ram.memory\[41\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05199__A2 _01777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09751_ _00145_ io_in[4] u_cpu.rf_ram.memory\[7\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06963_ _03110_ _03127_ _03133_ _00410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08137__A2 _02915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08702_ u_arbiter.i_wb_cpu_dbus_adr\[8\] u_arbiter.i_wb_cpu_dbus_adr\[9\] _04257_
+ _04264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05914_ _02443_ _00049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09682_ u_cpu.rf_ram.memory\[23\]\[4\] _04832_ _04837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06894_ u_cpu.rf_ram.memory\[64\]\[2\] _03089_ _03092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08633_ _03922_ _04188_ _04221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05845_ _02403_ u_cpu.cpu.genblk3.csr.i_mtip _02404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06699__A2 _02978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07896__A1 _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08564_ _02392_ _02320_ _03896_ _04161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05776_ _02347_ _02350_ _02351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_54_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07515_ _03322_ _03435_ _03443_ _00652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08696__I0 u_arbiter.i_wb_cpu_dbus_adr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08495_ _04096_ _04097_ _03966_ _04098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_23_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07446_ u_cpu.rf_ram.memory\[49\]\[0\] _03405_ _03406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06320__A1 _02657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07377_ _02637_ _03365_ _03367_ _00590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_136_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04882__A1 _01438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09116_ _04448_ _04503_ _04510_ _01187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06328_ u_cpu.rf_ram.memory\[80\]\[0\] _02756_ _02757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07820__A1 _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06623__A2 _02935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09047_ u_arbiter.i_wb_cpu_ibus_adr\[1\] u_arbiter.i_wb_cpu_ack _02461_ _04473_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_11_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06259_ u_cpu.rf_ram.memory\[18\]\[6\] _02707_ _02714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10747__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09573__A1 _04630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08376__A2 _03972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06387__A1 _02693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09949_ _00343_ io_in[4] u_cpu.rf_ram.memory\[6\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08128__A2 _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05336__B _01519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06139__A1 _02608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10897__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09628__A2 _04802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10127__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09322__I _02636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07639__A1 _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08836__B1 _04329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08300__A2 u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10724_ _00021_ io_in[4] u_cpu.cpu.alu.add_cy_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10655_ _01028_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06862__A2 _03069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10277__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08382__B _04003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04873__A1 u_cpu.cpu.state.genblk1.misalign_trap_sync_r vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08064__A1 _03695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10586_ _00959_ io_in[4] u_cpu.cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06614__A2 _02754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09564__A1 _02677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11138_ _00071_ io_in[0] u_scanchain_local.module_data_in\[50\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09316__A1 _04450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08119__A2 _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11069_ u_cpu.rf_ram_if.wdata0_r\[6\] io_in[4] u_cpu.rf_ram_if.wdata0_r\[5\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07878__A1 _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05630_ _01492_ _02179_ _02188_ _02207_ _02208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_92_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06550__A1 _02887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11052__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05561_ _01490_ _02130_ _02139_ _02140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_07300_ _02768_ _02838_ _03324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05492_ _01492_ _02062_ _02071_ _02072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_20_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08280_ _02909_ u_arbiter.i_wb_cpu_rdt\[15\] _03907_ _03908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_32_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06302__A1 _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07231_ _03108_ _03277_ _03282_ _00529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09912__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07162_ u_cpu.rf_ram.memory\[52\]\[6\] _03237_ _03244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06113_ _02361_ _02601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07802__A1 _02291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07093_ _03114_ _03197_ _03205_ _00468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06044_ u_cpu.cpu.ctrl.o_ibus_adr\[22\] _02541_ _02544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08512__S _02466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09555__A1 _04630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08358__A2 _03956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09803_ _00197_ io_in[4] u_cpu.rf_ram.memory\[44\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_101_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07030__A2 _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07995_ u_cpu.rf_ram.memory\[121\]\[3\] _03720_ _03724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__04919__A2 u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05041__A1 _01617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09734_ _00128_ io_in[4] u_cpu.rf_ram.memory\[20\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05156__B _01481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06946_ u_cpu.rf_ram.memory\[63\]\[6\] _03117_ _03124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09665_ _04632_ _04822_ _04827_ _01419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07869__A1 u_cpu.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06877_ _02887_ _03079_ _03082_ _00375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__04995__B _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08616_ _04203_ _04205_ _04206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_27_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05828_ io_in[3] _02388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09596_ u_cpu.rf_ram.memory\[24\]\[6\] _04782_ _04789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06541__A1 _02619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08547_ _02320_ _04144_ _04145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08818__B1 _04329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05759_ u_cpu.cpu.state.o_cnt_r\[0\] _02292_ _02334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08294__A1 _02464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07097__A2 _03207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08478_ _03912_ _04075_ _04082_ _03896_ _04083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_11_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07429_ _03306_ _03395_ _03396_ _00613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06844__A2 _03059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08046__A1 _03695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10440_ _00813_ io_in[4] u_cpu.rf_ram.memory\[35\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08597__A2 _03985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10371_ _00744_ io_in[4] u_cpu.rf_ram.memory\[123\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05280__A1 _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09546__A1 _02677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08349__A2 u_arbiter.i_wb_cpu_rdt\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09317__I _02631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07021__A2 _03157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05583__A2 _02161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11075__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08377__B _03998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05513__C _01486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09935__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08285__A1 _02465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07088__A2 _03197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05099__A1 _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10707_ _01077_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10912__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10638_ _01011_ io_in[4] u_cpu.rf_ram.memory\[31\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09085__I0 u_arbiter.i_wb_cpu_rdt\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04924__I _01499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04941__S1 _01525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08588__A2 _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10569_ _00942_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06599__A1 _01441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07260__A2 _03297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05271__A1 _01566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09537__A1 _04630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07012__A2 _03157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05023__A1 _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06800_ u_cpu.rf_ram.memory\[6\]\[0\] _03039_ _03040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07780_ u_cpu.rf_ram.memory\[36\]\[1\] _03593_ _03595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05574__A2 _02152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04992_ _01498_ _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06731_ u_cpu.rf_ram.memory\[77\]\[2\] _02998_ _03001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09450_ _04638_ _04691_ _04699_ _01332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06662_ _02891_ _02956_ _02961_ _00281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10442__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08401_ u_arbiter.i_wb_cpu_rdt\[21\] u_arbiter.i_wb_cpu_rdt\[5\] _02467_ _04020_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_24_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05613_ u_cpu.rf_ram.memory\[32\]\[7\] u_cpu.rf_ram.memory\[33\]\[7\] u_cpu.rf_ram.memory\[34\]\[7\]
+ u_cpu.rf_ram.memory\[35\]\[7\] _01495_ _01499_ _02191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09381_ u_cpu.rf_ram.memory\[85\]\[0\] _04661_ _04662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06593_ u_arbiter.i_wb_cpu_dbus_dat\[4\] _02916_ _02917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08332_ _02909_ u_arbiter.i_wb_cpu_rdt\[4\] _03957_ _03958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05544_ _01512_ _02122_ _02123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08276__A1 _03901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07079__A2 _03197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10592__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08263_ _03705_ _03885_ _03892_ _00952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05629__A3 _02206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06826__A2 _03049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05475_ _01464_ _02054_ _02055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07214_ u_cpu.rf_ram.memory\[142\]\[5\] _03267_ _03273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08028__A1 _02637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08194_ _03848_ _03849_ _00926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08579__A2 _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07145_ _03112_ _03227_ _03234_ _00491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05866__S _02418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07251__A2 _03287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07076_ _02827_ _02954_ _03196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05262__A1 _01548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09528__A1 _02677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06027_ _02528_ _02521_ _02529_ _02530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09808__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07003__A2 _03147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11098__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07978_ _03699_ _03710_ _03714_ _00845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09073__S _04485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09717_ _00111_ io_in[4] u_cpu.rf_ram.memory\[21\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06929_ _02666_ _03114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09958__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09700__A1 _02912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09648_ u_cpu.rf_ram.memory\[100\]\[5\] _04812_ _04818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05614__B _01518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06514__A1 _02687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10935__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09579_ _04636_ _04772_ _04779_ _01381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08644__C _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05876__I0 u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07490__A2 _03425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10423_ _00796_ io_in[4] u_cpu.rf_ram.memory\[90\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10354_ _00740_ io_in[4] u_cpu.rf_ram.memory\[124\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07242__A2 _03287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10315__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09519__A1 _01477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05253__A1 _01528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08990__A2 _04436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10285_ _00671_ io_in[4] u_cpu.rf_ram.memory\[131\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05005__A1 _01512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10465__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06808__A2 _03039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05260_ _01543_ _01841_ _01842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05492__A1 _01492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05191_ u_cpu.rf_ram.memory\[100\]\[2\] u_cpu.rf_ram.memory\[101\]\[2\] u_cpu.rf_ram.memory\[102\]\[2\]
+ u_cpu.rf_ram.memory\[103\]\[2\] _01551_ _01573_ _01774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08570__B _04165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07233__A2 _03277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08430__A1 _03697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05244__A1 _01506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08981__A2 _04425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08950_ u_cpu.cpu.immdec.imm11_7\[3\] _04390_ _04411_ _03955_ _04412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__10808__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07901_ u_cpu.rf_ram.memory\[35\]\[5\] _03662_ _03668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08881_ _02647_ _04361_ _04365_ _01097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07832_ _03510_ _03616_ _03624_ _00788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07763_ _03498_ _03583_ _03585_ _00758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10958__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04975_ _01540_ _01560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09502_ _04732_ _02303_ _01458_ _02305_ _04733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_25_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06714_ _02887_ _02988_ _02991_ _00303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08497__A1 _01444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07694_ u_cpu.rf_ram.memory\[125\]\[3\] _03543_ _03547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09433_ _02870_ _04349_ _04690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06645_ _02893_ _02945_ _02951_ _00274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09364_ _02632_ _04651_ _04652_ _01293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_75_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06576_ u_cpu.rf_ram.memory\[4\]\[4\] _02900_ _02905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08315_ _02465_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[3\] _03943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05527_ u_cpu.rf_ram.memory\[40\]\[6\] u_cpu.rf_ram.memory\[41\]\[6\] u_cpu.rf_ram.memory\[42\]\[6\]
+ u_cpu.rf_ram.memory\[43\]\[6\] _01551_ _01524_ _02106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09295_ u_cpu.rf_ram.memory\[108\]\[6\] _04603_ _04610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08246_ u_arbiter.i_wb_cpu_rdt\[31\] _02924_ _03874_ _02277_ _03883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_36_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05458_ _01548_ _02037_ _01579_ _02038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_20_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07472__A2 _03415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10338__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08177_ u_arbiter.i_wb_cpu_dbus_dat\[7\] _03835_ _03838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05389_ _01597_ _01969_ _01600_ _01970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_21_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07128_ u_cpu.rf_ram.memory\[54\]\[7\] _03217_ _03225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08421__A1 _03965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07224__A2 _03277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05235__A1 _01465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08972__A2 _04425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05609__B _01481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07059_ _03186_ _03187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10488__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05786__A2 u_cpu.cpu.ctrl.i_iscomp vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06983__A1 _03112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10070_ _00464_ io_in[4] u_cpu.rf_ram.memory\[56\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08700__S _04257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09780__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05094__S0 _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10972_ _01341_ io_in[4] u_cpu.rf_ram.memory\[88\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08488__A1 u_cpu.cpu.immdec.imm24_20\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08488__B2 u_cpu.cpu.immdec.imm30_25\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05397__S1 _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11113__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08660__A1 _03699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10406_ _00779_ io_in[4] u_cpu.cpu.state.o_cnt_r\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07215__A2 _03267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05226__A1 _01512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10337_ _00723_ io_in[4] u_cpu.rf_ram.memory\[126\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08963__A2 _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05777__A2 _02305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10268_ _00654_ io_in[4] u_cpu.rf_ram.memory\[133\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05238__C _01466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10199_ _00585_ io_in[4] u_cpu.rf_ram.memory\[143\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05085__S0 _01495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08479__A1 u_cpu.cpu.immdec.imm24_20\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09140__A2 _04523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05388__S1 _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07151__A1 _03098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06430_ u_cpu.rf_ram.memory\[44\]\[1\] _02816_ _02818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05701__A2 _02277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06361_ _02689_ _02770_ _02776_ _00165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08100_ _03695_ _03780_ _03782_ _00899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05312_ _01621_ _01893_ _01894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09080_ _04491_ _01170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07454__A2 _03405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06292_ _02637_ _02733_ _02735_ _00137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08651__A1 _02754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05465__A1 _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08031_ u_cpu.rf_ram.memory\[11\]\[3\] _03740_ _03744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05243_ u_cpu.rf_ram.memory\[24\]\[3\] u_cpu.rf_ram.memory\[25\]\[3\] u_cpu.rf_ram.memory\[26\]\[3\]
+ u_cpu.rf_ram.memory\[27\]\[3\] _01508_ _01509_ _01825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10630__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08403__A1 _04000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07206__A2 _03267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05174_ _01548_ _01756_ _01518_ _01757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_115_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05217__A1 _01617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08954__A2 _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09982_ _00376_ io_in[4] u_cpu.rf_ram.memory\[65\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05429__B _01534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06965__A1 _03112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08933_ _03910_ _04395_ _03965_ _04396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__04976__B1 _01553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10780__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08167__B1 _03808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08864_ u_cpu.rf_ram.memory\[109\]\[4\] _04351_ _04356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05076__S0 _01530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07815_ _02626_ _02849_ _03615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08795_ _04317_ _01059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__07390__A1 _02780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10010__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11136__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07746_ u_cpu.rf_ram.memory\[38\]\[2\] _03573_ _03576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04958_ _01463_ _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09131__A2 _04513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07677_ _03502_ _03533_ _03537_ _00720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_77_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_04889_ u_cpu.cpu.decode.op26 u_cpu.cpu.decode.co_ebreak _01476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09416_ _04680_ _04681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06628_ u_cpu.rf_ram.memory\[16\]\[6\] _02935_ _02942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07693__A2 _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08890__A1 _02619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10160__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09347_ u_cpu.rf_ram.memory\[59\]\[1\] _04641_ _04643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06559_ _02893_ _02883_ _02894_ _00245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08642__A1 _04165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09278_ _04448_ _04593_ _04600_ _01259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05456__A1 _01512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05000__S0 _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08229_ u_arbiter.i_wb_cpu_rdt\[24\] _03807_ _03808_ u_arbiter.i_wb_cpu_dbus_dat\[24\]
+ _03873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_5_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09198__A2 _04553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05759__A2 _02292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10122_ _00516_ io_in[4] u_cpu.rf_ram.memory\[15\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10053_ _00447_ io_in[4] u_cpu.rf_ram.memory\[58\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09325__I _02641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05067__S0 _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09370__A2 _04651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07381__A1 _02647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06184__A2 _02628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05931__A2 _02403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09122__A2 _04513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10955_ _01324_ io_in[4] u_cpu.rf_ram.memory\[86\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10503__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07133__A1 _03098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07684__A2 _03533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08881__A1 _02647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10886_ _01255_ io_in[4] u_cpu.rf_ram.memory\[83\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10653__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08633__A1 _03922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07436__A2 _03395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08484__I1 u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05447__A1 _01548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05998__A2 _02499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09189__A2 _04543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11009__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06947__A1 _03112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05930_ _02403_ u_scanchain_local.module_data_in\[36\] _02453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10033__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05058__S0 _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09361__A2 _02780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05861_ _02414_ _02403_ _02408_ _02415_ _00081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07372__A1 _02731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07600_ u_cpu.rf_ram.memory\[12\]\[5\] _03485_ _03491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_94_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08580_ _04171_ _04165_ _04172_ _04008_ _00989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05792_ _00798_ _02358_ _02365_ _02366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09113__A2 _04503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07531_ _03320_ _03445_ _03452_ _00659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10183__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05712__B _02286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07462_ _02954_ _02976_ _03414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07675__A2 _03533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08872__A1 _02731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09201_ u_cpu.rf_ram.memory\[79\]\[4\] _04553_ _04558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06413_ u_cpu.rf_ram.memory\[45\]\[2\] _02805_ _02808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05230__S0 _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07393_ _03306_ _03375_ _03376_ _00597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09132_ _04446_ _04513_ _04519_ _01194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05781__S1 _02355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06344_ _02609_ _02613_ _02765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08624__A1 _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05438__A1 _01504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09063_ _04446_ _04476_ _04482_ _01162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06275_ u_cpu.rf_ram.memory\[20\]\[4\] _02719_ _02724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08014_ _02647_ _03730_ _03734_ _00861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_135_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05226_ _01512_ _01808_ _01481_ _01809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05157_ u_cpu.rf_ram.memory\[20\]\[2\] u_cpu.rf_ram.memory\[21\]\[2\] u_cpu.rf_ram.memory\[22\]\[2\]
+ u_cpu.rf_ram.memory\[23\]\[2\] _01497_ _01501_ _01740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_89_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05874__S _02418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09965_ _00359_ io_in[4] u_cpu.rf_ram.memory\[67\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05088_ _01505_ _01671_ _01672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08916_ u_cpu.rf_ram.memory\[93\]\[3\] _04381_ _04385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09896_ _00290_ io_in[4] u_cpu.rf_ram.memory\[119\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09352__A2 _04641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10526__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08847_ _04344_ _01084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__07363__A1 _03314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06166__A2 _02628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08560__B1 _03909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08778_ u_cpu.rf_ram.memory\[30\]\[7\] _04299_ _04307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09081__S _04485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09104__A2 _04503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07729_ _03500_ _03563_ _03566_ _00743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07115__A1 _03098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10676__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10740_ _01109_ io_in[4] u_cpu.rf_ram.memory\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08863__A1 _03699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07666__A2 _03523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05516__I2 u_cpu.rf_ram.memory\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05677__A1 _01465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05221__S0 _01507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10671_ _00022_ io_in[4] u_cpu.cpu.bufreg.c_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08933__B _03965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08615__A1 _04031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07418__A2 _03385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05429__A1 _01528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08091__A2 _03770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08918__A2 _04381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10056__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09040__A1 _04446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05288__S0 _01496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09591__A2 _04782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08394__A3 _04013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11154_ _00088_ io_in[0] u_scanchain_local.module_data_in\[66\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10105_ _00499_ io_in[4] u_cpu.rf_ram.memory\[52\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11085_ u_cpu.cpu.o_wen0 io_in[4] u_cpu.rf_ram_if.wen0_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10036_ _00430_ io_in[4] u_cpu.rf_ram.memory\[19\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09343__A2 _02849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07354__A1 _02870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04927__I _01463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10938_ _01307_ io_in[4] u_cpu.rf_ram.memory\[85\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08854__A1 _02803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07657__A2 _03523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05668__A1 _01492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05212__S0 _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10869_ _01238_ io_in[4] u_cpu.rf_ram.memory\[106\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08606__A1 _03912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04891__A2 _01477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08082__A2 _03770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06093__A1 _02463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06060_ _02553_ _02557_ _00084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_126_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05011_ _01543_ _01595_ _01596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05279__S0 _01551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09582__A2 _02954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10549__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06396__A2 _02794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07593__A1 _02637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08790__B1 _04311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09750_ _00144_ io_in[4] u_cpu.rf_ram.memory\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06962_ u_cpu.rf_ram.memory\[62\]\[5\] _03127_ _03133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09841__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05913_ u_arbiter.i_wb_cpu_rdt\[27\] u_arbiter.i_wb_cpu_dbus_dat\[24\] _02431_ _02443_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08701_ _04263_ _01019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09681_ _04630_ _04832_ _04836_ _01426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06893_ _02885_ _03089_ _03091_ _00382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06148__A2 _02628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07345__A1 _03314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08632_ _04165_ _04218_ _04219_ _04220_ _00993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_66_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10699__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05844_ _02402_ _02403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07896__A2 _03662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08563_ _03925_ _04009_ _04158_ _04159_ _04160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05775_ _01443_ _02348_ _02349_ _02334_ _02336_ _02350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_70_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09991__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07514_ u_cpu.rf_ram.memory\[134\]\[7\] _03435_ _03443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05442__B _01558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08494_ _03935_ _03914_ _03903_ _03961_ _04097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07648__A2 _03513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07445_ _03404_ _03405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05161__C _01486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06320__A2 _02745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07376_ u_cpu.rf_ram.memory\[14\]\[1\] _03365_ _03367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09115_ u_cpu.rf_ram.memory\[101\]\[6\] _04503_ _04510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04882__A2 _01452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06327_ _02755_ _02756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10079__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08073__A2 _03760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09270__A1 _04440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06084__A1 _02389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09046_ _04141_ _04472_ _01155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06258_ _02689_ _02707_ _02713_ _00125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07820__A2 _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05209_ _01490_ _01782_ _01791_ _01792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05831__A1 _01441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09022__A1 _04446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05831__B2 _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06189_ _02666_ _02667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09573__A2 _04772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06387__A2 _02784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09948_ _00342_ io_in[4] u_cpu.rf_ram.memory\[6\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09879_ _00273_ io_in[4] u_cpu.rf_ram.memory\[17\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07336__A1 _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07887__A2 _03652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07639__A2 _03513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10723_ _01093_ io_in[4] u_cpu.rf_ram.memory\[109\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06311__A2 _02745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10654_ _01027_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09714__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08064__A2 _03760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10585_ _00958_ io_in[4] u_cpu.cpu.branch_op vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06075__A1 _02403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09864__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09564__A2 _02838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06378__A2 _02784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07575__A1 _03310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11137_ _00069_ io_in[0] u_scanchain_local.module_data_in\[49\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10841__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09316__A2 _04613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11068_ u_cpu.rf_ram_if.wdata0_r\[5\] io_in[4] u_cpu.rf_ram_if.wdata0_r\[4\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07327__A1 _03314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10019_ _00413_ io_in[4] u_cpu.rf_ram.memory\[61\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07878__A2 _03652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10991__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06550__A2 _02883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05262__B _01518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05560_ _02132_ _02134_ _02136_ _02138_ _01581_ _02139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_17_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05491_ _02064_ _02066_ _02068_ _02070_ _01541_ _02071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_60_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06302__A2 _02733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08573__B _04165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07230_ u_cpu.rf_ram.memory\[141\]\[4\] _03277_ _03282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10221__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07161_ _03110_ _03237_ _03243_ _00498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09252__A1 _04440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08055__A2 _03750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06112_ u_cpu.cpu.ctrl.pc_plus_4_cy_r u_arbiter.i_wb_cpu_ibus_adr\[0\] _02600_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07092_ u_cpu.rf_ram.memory\[56\]\[7\] _03197_ _03205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07802__A2 _03605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10371__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05813__A1 _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06043_ _02540_ _02542_ _02543_ _00080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09555__A2 _04762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09802_ _00196_ io_in[4] u_cpu.rf_ram.memory\[44\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07994_ _03697_ _03720_ _03723_ _00852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09307__A2 _04613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05672__S0 _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06945_ _03110_ _03117_ _03123_ _00402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09733_ _00127_ io_in[4] u_cpu.rf_ram.memory\[18\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07318__A1 _02743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08748__B _02598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09664_ u_cpu.rf_ram.memory\[89\]\[4\] _04822_ _04827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06876_ u_cpu.rf_ram.memory\[65\]\[2\] _03079_ _03082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07869__A2 _03611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08615_ _04031_ _04204_ _04205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05827_ _01467_ _02379_ _02387_ _00014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09595_ _04634_ _04782_ _04788_ _01388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06541__A2 _02827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08546_ _01444_ _02265_ u_cpu.cpu.decode.opcode\[1\] _04144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05758_ _02317_ _02319_ _02324_ _02332_ _02333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_35_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09737__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08477_ _04031_ _04078_ _04080_ _04081_ _03912_ _04082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_05689_ _01444_ _02265_ u_cpu.cpu.decode.opcode\[1\] _02266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_126_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07428_ u_cpu.rf_ram.memory\[137\]\[0\] _03395_ _03396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10714__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07359_ _03310_ _03355_ _03357_ _00582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08046__A2 _03750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09887__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10370_ _00743_ io_in[4] u_cpu.rf_ram.memory\[123\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09029_ u_cpu.rf_ram.memory\[96\]\[0\] _04463_ _04464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05804__A1 _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10864__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09546__A2 _02780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07557__A1 _03310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05663__S0 _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07309__A1 _03314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08377__C _03922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06532__A2 _02872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10244__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09482__A1 _04634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06296__A1 _02647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10706_ _01076_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10394__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09234__A1 _04440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10637_ _01010_ io_in[4] u_cpu.rf_ram.memory\[31\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08037__A2 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10568_ _00941_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06599__A2 _02309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10499_ _00872_ io_in[4] u_cpu.rf_ram.memory\[11\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09537__A2 _04752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04940__I _01524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05257__B _01482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05023__A2 _01606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05654__S0 _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_04991_ _01495_ _01576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_49_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06771__A2 _03018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08568__B _02911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06730_ _02885_ _02998_ _03000_ _00310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_49_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05406__S0 _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06661_ u_cpu.rf_ram.memory\[40\]\[4\] _02956_ _02961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08400_ _02325_ _03956_ _04019_ _00962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05612_ _01571_ _02189_ _02190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09380_ _04660_ _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_91_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06592_ u_arbiter.i_wb_cpu_dbus_dat\[3\] u_arbiter.i_wb_cpu_dbus_dat\[2\] u_arbiter.i_wb_cpu_dbus_dat\[0\]
+ u_arbiter.i_wb_cpu_dbus_dat\[1\] _02916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_24_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05582__I0 u_cpu.rf_ram.memory\[128\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08331_ _02466_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[4\] _03957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_51_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05543_ u_cpu.rf_ram.memory\[100\]\[6\] u_cpu.rf_ram.memory\[101\]\[6\] u_cpu.rf_ram.memory\[102\]\[6\]
+ u_cpu.rf_ram.memory\[103\]\[6\] _01551_ _01524_ _02122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10737__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08276__A2 _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06287__A1 _02695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08262_ u_cpu.rf_ram.memory\[113\]\[6\] _03885_ _03892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05720__B _02292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05474_ u_cpu.rf_ram.memory\[92\]\[5\] u_cpu.rf_ram.memory\[93\]\[5\] u_cpu.rf_ram.memory\[94\]\[5\]
+ u_cpu.rf_ram.memory\[95\]\[5\] _01562_ _01563_ _02054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07213_ _03108_ _03267_ _03272_ _00521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08193_ u_arbiter.i_wb_cpu_rdt\[12\] _03822_ _03833_ u_arbiter.i_wb_cpu_dbus_dat\[13\]
+ _03849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08028__A2 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07144_ u_cpu.rf_ram.memory\[53\]\[6\] _03227_ _03234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10887__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07787__A1 _03504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07075_ _03114_ _03187_ _03195_ _00460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05946__I _02465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09528__A2 _02849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05262__A2 _01843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06026_ u_cpu.cpu.ctrl.o_ibus_adr\[19\] _02529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_126_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10117__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07539__A1 _03310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05882__S _02418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07977_ u_cpu.rf_ram.memory\[118\]\[3\] _03710_ _03714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09716_ _00110_ io_in[4] u_cpu.rf_ram.memory\[21\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10267__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06928_ _03112_ _03100_ _03113_ _00395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05970__B1 _02398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09647_ _04632_ _04812_ _04817_ _01411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_16_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06859_ _02887_ _03069_ _03072_ _00367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_16_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07711__A1 _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06514__A2 _02861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09578_ u_cpu.rf_ram.memory\[25\]\[6\] _04772_ _04779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08529_ _03935_ _03974_ _04052_ _04128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09464__A1 _04634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08267__A2 _02461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06278__A1 _02689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05630__B _02207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05876__I1 u_arbiter.i_wb_cpu_dbus_dat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08019__A2 _03730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09216__A1 _04440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08941__B _03965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10422_ _00795_ io_in[4] u_cpu.rf_ram.memory\[90\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10353_ _00739_ io_in[4] u_cpu.rf_ram.memory\[124\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05856__I _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09328__I _02646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05253__A2 _01834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06450__A1 _02669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10284_ _00670_ io_in[4] u_cpu.rf_ram.memory\[131\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11042__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05077__B _01534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05005__A2 _01589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07950__A1 _03695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08388__B _04008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06753__A2 _03008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09902__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06505__A2 _02861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05159__I3 u_cpu.rf_ram.memory\[19\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08258__A2 _03885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05190_ _01492_ _01744_ _01753_ _01772_ _01773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_127_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07769__A1 _03504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08430__A2 _04041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05244__A2 _01825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06441__A1 _02691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06992__A2 _03147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07900_ _03504_ _03662_ _03667_ _00814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08880_ u_cpu.rf_ram.memory\[3\]\[3\] _04361_ _04365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07831_ u_cpu.rf_ram.memory\[91\]\[7\] _03616_ _03624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04974_ _01554_ _01557_ _01558_ _01559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07762_ u_cpu.rf_ram.memory\[37\]\[1\] _03583_ _03585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09501_ u_cpu.cpu.genblk3.csr.mcause3_0\[3\] _04732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06713_ u_cpu.rf_ram.memory\[139\]\[2\] _02988_ _02991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07693_ _03500_ _03543_ _03546_ _00727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05434__C _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08497__A2 _02305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09432_ _04638_ _04681_ _04689_ _01324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06644_ u_cpu.rf_ram.memory\[17\]\[5\] _02945_ _02951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06575_ _02647_ _02900_ _02904_ _00251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_24_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09363_ u_cpu.rf_ram.memory\[10\]\[0\] _04651_ _04652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09446__A1 _04634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08314_ _03940_ _03941_ _03942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_05526_ _01504_ _02104_ _01518_ _02105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09294_ _04446_ _04603_ _04609_ _01266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08245_ _02450_ _03835_ _03833_ _02452_ _03882_ _00944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_05457_ u_cpu.rf_ram.memory\[96\]\[5\] u_cpu.rf_ram.memory\[97\]\[5\] u_cpu.rf_ram.memory\[98\]\[5\]
+ u_cpu.rf_ram.memory\[99\]\[5\] _01567_ _01568_ _02037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_21_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05322__I3 u_cpu.rf_ram.memory\[139\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06680__A1 u_cpu.rf_ram.memory\[119\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08176_ _03836_ _03837_ _00920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05388_ u_cpu.rf_ram.memory\[88\]\[4\] u_cpu.rf_ram.memory\[89\]\[4\] u_cpu.rf_ram.memory\[90\]\[4\]
+ u_cpu.rf_ram.memory\[91\]\[4\] _01598_ _01556_ _01969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_10_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11065__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07127_ _03112_ _03217_ _03224_ _00483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08421__A2 _04030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05235__A2 _01817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07058_ _02827_ _02838_ _03186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06009_ u_cpu.cpu.ctrl.o_ibus_adr\[15\] u_cpu.cpu.ctrl.o_ibus_adr\[14\] _02508_ _02515_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06983__A2 _03137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09925__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06735__A2 _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07932__A1 _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10902__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05094__S1 _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10971_ _01340_ io_in[4] u_cpu.rf_ram.memory\[87\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09685__A1 _04634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08488__A2 _04069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07160__A2 _03237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08660__A2 _04237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10405_ _00778_ io_in[4] u_cpu.cpu.state.o_cnt_r\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10432__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05226__A2 _01808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10336_ _00722_ io_in[4] u_cpu.rf_ram.memory\[126\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05777__A3 _02265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06974__A2 _03137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10267_ _00653_ io_in[4] u_cpu.rf_ram.memory\[133\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04985__A1 _01566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10582__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10198_ _00584_ io_in[4] u_cpu.rf_ram.memory\[143\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05535__B _01480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05085__S1 _01499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08479__A2 _03955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07151__A2 _03237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09428__A1 _04634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06360_ u_cpu.rf_ram.memory\[78\]\[5\] _02770_ _02776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08100__A1 _03695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11088__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05311_ u_cpu.rf_ram.memory\[72\]\[3\] u_cpu.rf_ram.memory\[73\]\[3\] u_cpu.rf_ram.memory\[74\]\[3\]
+ u_cpu.rf_ram.memory\[75\]\[3\] _01562_ _01622_ _01893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_30_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06291_ u_cpu.rf_ram.memory\[1\]\[1\] _02733_ _02735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08651__A2 _02782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08030_ _02642_ _03740_ _03743_ _00868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05465__A2 _02044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05242_ _01493_ _01823_ _01824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06662__A1 _02891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09948__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05173_ u_cpu.rf_ram.memory\[32\]\[2\] u_cpu.rf_ram.memory\[33\]\[2\] u_cpu.rf_ram.memory\[34\]\[2\]
+ u_cpu.rf_ram.memory\[35\]\[2\] _01495_ _01499_ _01756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09600__A1 _02731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05217__A2 _01799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06414__A1 _02683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09981_ _00375_ io_in[4] u_cpu.rf_ram.memory\[65\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06965__A2 _03127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10925__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08932_ _03928_ _04188_ _04190_ _04394_ _03969_ _04395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_88_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08167__A1 u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08167__B2 u_arbiter.i_wb_cpu_dbus_dat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08863_ _03699_ _04351_ _04355_ _01089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06717__A2 _02988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07914__A1 _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07814_ _03614_ _00780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05076__S1 _01532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08794_ u_cpu.cpu.ctrl.o_ibus_adr\[5\] _04309_ _04311_ u_cpu.cpu.ctrl.o_ibus_adr\[6\]
+ _04317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07390__A2 _02976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04957_ _01527_ _01535_ _01537_ _01539_ _01541_ _01542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_42_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07745_ _03498_ _03573_ _03575_ _00750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09667__A1 _04634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08714__I0 u_arbiter.i_wb_cpu_dbus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07676_ u_cpu.rf_ram.memory\[126\]\[3\] _03533_ _03537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04888_ u_cpu.cpu.immdec.imm24_20\[1\] _01475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07142__A2 _03227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09415_ _02626_ _03037_ _04680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10305__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06627_ _02893_ _02935_ _02941_ _00266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08890__A2 _02731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06558_ u_cpu.rf_ram.memory\[50\]\[5\] _02883_ _02894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09346_ _04622_ _04641_ _04642_ _01285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05509_ u_cpu.rf_ram.memory\[20\]\[6\] u_cpu.rf_ram.memory\[21\]\[6\] u_cpu.rf_ram.memory\[22\]\[6\]
+ u_cpu.rf_ram.memory\[23\]\[6\] _01530_ _01501_ _02088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09277_ u_cpu.rf_ram.memory\[83\]\[6\] _04593_ _04600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06489_ u_cpu.rf_ram.memory\[43\]\[1\] _02851_ _02853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08491__B _03899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10455__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09079__S _04485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05000__S1 _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08228_ u_arbiter.i_wb_cpu_dbus_dat\[25\] _03833_ _03872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08159_ _02915_ _02916_ _03823_ _03824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_134_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06405__A1 _02693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10121_ _00515_ io_in[4] u_cpu.rf_ram.memory\[15\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06956__A2 _03127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08158__A1 u_arbiter.i_wb_cpu_dbus_dat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10052_ _00446_ io_in[4] u_cpu.rf_ram.memory\[58\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05067__S1 _01509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07381__A2 _03365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10954_ _01323_ io_in[4] u_cpu.rf_ram.memory\[86\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07133__A2 _03227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08881__A2 _04361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10885_ _01254_ io_in[4] u_cpu.rf_ram.memory\[83\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05090__B _01558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10948__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08397__A1 _02911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06205__I _02636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05249__C _01486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06947__A2 _03117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10319_ _00705_ io_in[4] u_cpu.rf_ram.memory\[128\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05860_ u_cpu.cpu.bne_or_bge _02306_ _02355_ _02415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05058__S1 _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07372__A2 _02766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10328__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09649__A1 _04634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05383__A1 _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05791_ _02363_ _02364_ _01460_ _02300_ _02365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_81_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08576__B _04165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07530_ u_cpu.rf_ram.memory\[133\]\[6\] _03445_ _03452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08321__A1 _03906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07124__A2 _03217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07461_ _03322_ _03405_ _03413_ _00628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08872__A2 _02825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09200_ _04442_ _04553_ _04557_ _01224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10478__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06412_ _02681_ _02805_ _02807_ _00185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_16_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06883__A1 _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07392_ u_cpu.rf_ram.memory\[138\]\[0\] _03375_ _03376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05230__S1 _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09131_ u_cpu.rf_ram.memory\[102\]\[5\] _04513_ _04519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06343_ _02693_ _02756_ _02764_ _00159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09770__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08624__A2 _03975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09062_ u_cpu.rf_ram.memory\[28\]\[5\] _04476_ _04482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06635__A1 _02881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05438__A2 _02017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06274_ _02685_ _02719_ _02723_ _00131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05225_ u_cpu.rf_ram.memory\[76\]\[2\] u_cpu.rf_ram.memory\[77\]\[2\] u_cpu.rf_ram.memory\[78\]\[2\]
+ u_cpu.rf_ram.memory\[79\]\[2\] _01529_ _01500_ _01808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08013_ u_cpu.rf_ram.memory\[8\]\[3\] _03730_ _03734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08388__A1 _02309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05156_ _01506_ _01738_ _01481_ _01739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06938__A2 _03117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09964_ _00358_ io_in[4] u_cpu.rf_ram.memory\[67\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05087_ u_cpu.rf_ram.memory\[40\]\[1\] u_cpu.rf_ram.memory\[41\]\[1\] u_cpu.rf_ram.memory\[42\]\[1\]
+ u_cpu.rf_ram.memory\[43\]\[1\] _01551_ _01524_ _01671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__11103__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08915_ _03697_ _04381_ _04384_ _01112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08330__I _03955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09895_ _00289_ io_in[4] u_cpu.rf_ram.memory\[119\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08846_ u_cpu.cpu.ctrl.o_ibus_adr\[30\] _04327_ _04329_ u_cpu.cpu.ctrl.o_ibus_adr\[31\]
+ _04344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08560__A1 _03899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07363__A2 _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08560__B2 _03925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05374__A1 _01566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08777_ _03705_ _04299_ _04306_ _01052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05989_ u_cpu.cpu.ctrl.o_ibus_adr\[10\] _02493_ u_cpu.cpu.ctrl.o_ibus_adr\[11\] _02500_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_73_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08486__B _03938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07728_ u_cpu.rf_ram.memory\[123\]\[2\] _03563_ _03566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07115__A2 _03217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07659_ _03502_ _03523_ _03527_ _00712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08863__A2 _04351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05221__S1 _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10670_ _01043_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08706__S _04257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09329_ u_cpu.rf_ram.memory\[84\]\[3\] _04624_ _04631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05429__A2 _02008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08379__A1 _04000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08379__B2 _03944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08441__S _02466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09040__A2 _04463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07051__A1 _03108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05288__S1 _01594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11153_ _00087_ io_in[0] u_scanchain_local.module_data_in\[65\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10104_ _00498_ io_in[4] u_cpu.rf_ram.memory\[52\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11084_ u_cpu.cpu.o_wdata1 io_in[4] u_cpu.rf_ram_if.wdata1_r\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10035_ _00429_ io_in[4] u_cpu.rf_ram.memory\[19\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08551__A1 _03925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07354__A2 _02976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05365__A1 _01490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10620__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08303__A1 _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07106__A2 _03207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05117__A1 _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10937_ _01306_ io_in[4] u_cpu.rf_ram.memory\[85\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08854__A2 _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09793__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05212__S1 _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06865__A1 _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10868_ _01237_ io_in[4] u_cpu.rf_ram.memory\[106\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10770__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10799_ _01168_ io_in[4] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06617__A1 _02881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04943__I _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07290__A1 _03316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10000__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11126__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05010_ u_cpu.rf_ram.memory\[124\]\[0\] u_cpu.rf_ram.memory\[125\]\[0\] u_cpu.rf_ram.memory\[126\]\[0\]
+ u_cpu.rf_ram.memory\[127\]\[0\] _01496_ _01594_ _01595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_126_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09031__A2 _04463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05279__S1 _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07593__A2 _03485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10150__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06961_ _03108_ _03127_ _03132_ _00409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08700_ u_arbiter.i_wb_cpu_dbus_adr\[7\] u_arbiter.i_wb_cpu_dbus_adr\[8\] _04257_
+ _04263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05912_ _02442_ _00047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09680_ u_cpu.rf_ram.memory\[23\]\[3\] _04832_ _04836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06892_ u_cpu.rf_ram.memory\[64\]\[1\] _03089_ _03091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07345__A2 _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08631_ u_cpu.cpu.immdec.imm19_12_20\[7\] _04165_ _04220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05843_ _02401_ _02402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08562_ _03896_ _03912_ _04159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05774_ _01441_ _02309_ u_cpu.cpu.alu.cmp_r _02349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_35_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07513_ _03320_ _03435_ _03442_ _00651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05108__A1 _01512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08493_ _03901_ _04094_ _04095_ _04096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_126_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07444_ _02695_ _02827_ _03404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05903__I0 u_arbiter.i_wb_cpu_rdt\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07375_ _02632_ _03365_ _03366_ _00589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_31_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09114_ _04446_ _04503_ _04509_ _01186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06608__A1 _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04853__I u_cpu.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06326_ _02626_ _02754_ _02755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09270__A2 _04593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06257_ u_cpu.rf_ram.memory\[18\]\[5\] _02707_ _02713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09045_ u_cpu.cpu.bufreg.i_sh_signed _03897_ _04472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07281__A1 _03310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05208_ _01784_ _01786_ _01788_ _01790_ _01581_ _01791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_117_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05831__A2 _02355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06188_ _02665_ _02666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09022__A2 _04453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07033__A1 _02652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05139_ _01716_ _01718_ _01720_ _01722_ _01541_ _01723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_104_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07584__A2 _03475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09947_ _00341_ io_in[4] u_cpu.rf_ram.memory\[6\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09878_ _00272_ io_in[4] u_cpu.rf_ram.memory\[17\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10643__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08533__A1 _03908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07336__A2 _03037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08829_ _04335_ _01075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_85_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10793__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08836__A2 _04327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10722_ _01092_ io_in[4] u_cpu.rf_ram.memory\[109\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06847__A1 _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10653_ _01026_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__04953__S0 _01530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10023__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11149__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10584_ _00957_ io_in[4] u_arbiter.i_wb_cpu_dbus_we vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09261__A2 _04583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05822__A2 _01467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09013__A2 _04453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10173__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07575__A2 _03475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11136_ _00068_ io_in[0] u_scanchain_local.module_data_in\[48\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11067_ u_cpu.rf_ram_if.wdata0_r\[4\] io_in[4] u_cpu.rf_ram_if.wdata0_r\[3\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08524__A1 _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07327__A2 _03335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10018_ _00412_ io_in[4] u_cpu.rf_ram.memory\[62\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__04938__I _01522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05490_ _01617_ _02069_ _01481_ _02070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05197__S0 _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05510__A1 _01513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07160_ u_cpu.rf_ram.memory\[52\]\[5\] _03237_ _03243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09252__A2 _04583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10516__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06111_ _02597_ _02333_ _02599_ _00024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07263__A1 _02642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07091_ _03112_ _03197_ _03204_ _00467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06042_ _02402_ u_scanchain_local.module_data_in\[58\] _02478_ u_arbiter.i_wb_cpu_dbus_adr\[21\]
+ _02543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_126_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09004__A2 _04436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07015__A1 _03108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10666__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09801_ _00195_ io_in[4] u_cpu.rf_ram.memory\[44\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07566__A2 _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07993_ u_cpu.rf_ram.memory\[121\]\[2\] _03720_ _03723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09732_ _00126_ io_in[4] u_cpu.rf_ram.memory\[18\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05672__S1 _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06944_ u_cpu.rf_ram.memory\[63\]\[5\] _03117_ _03123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07318__A2 _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05009__I _01499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09663_ _04630_ _04822_ _04826_ _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06875_ _02885_ _03079_ _03081_ _00374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08614_ _04178_ _04180_ _03924_ _04204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_54_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05826_ u_cpu.rf_ram_if.rdata0\[7\] _01467_ _02387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09594_ u_cpu.rf_ram.memory\[24\]\[5\] _04782_ _04788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08545_ u_cpu.cpu.immdec.imm19_12_20\[0\] _04143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_36_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05757_ u_cpu.cpu.ctrl.pc_plus_offset_cy_r _02331_ _02332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_78_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08818__A2 _04327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10046__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06829__A1 _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08476_ _03941_ _04051_ _04075_ _03947_ _04031_ _04081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_126_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05688_ u_cpu.cpu.decode.opcode\[0\] _02265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07427_ _03394_ _03395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05501__A1 _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07358_ u_cpu.rf_ram.memory\[143\]\[1\] _03355_ _03357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09243__A2 _04573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10196__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06309_ u_cpu.rf_ram.memory\[7\]\[0\] _02745_ _02746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08451__B1 _03988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07289_ u_cpu.rf_ram.memory\[72\]\[4\] _03308_ _03317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09087__S _04485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09028_ _04462_ _04463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_3_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05804__A2 _02373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05360__S0 _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07557__A2 _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05112__S0 _01496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05663__S1 _01563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08506__A1 _04067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07309__A2 _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05363__B _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05082__C _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05740__A1 _01442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09482__A2 _04711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10539__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10705_ _01075_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06296__A2 _02733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07493__A1 _03318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10636_ _01009_ io_in[4] u_cpu.rf_ram.memory\[31\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09831__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09234__A2 _04573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07245__A1 _03104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10567_ _00940_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10689__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08993__A1 _04440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06599__A3 _02922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05351__S0 _01551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10498_ _00871_ io_in[4] u_cpu.rf_ram.memory\[11\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09981__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07548__A2 _03455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05103__S0 _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05559__A1 _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08849__B _01451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11119_ _00050_ io_in[0] u_arbiter.i_wb_cpu_rdt\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05654__S1 _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04990_ _01571_ _01574_ _01575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09170__A1 _04448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10069__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06660_ _02889_ _02956_ _02960_ _00280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05406__S1 _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07720__A2 _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05611_ u_cpu.rf_ram.memory\[36\]\[7\] u_cpu.rf_ram.memory\[37\]\[7\] u_cpu.rf_ram.memory\[38\]\[7\]
+ u_cpu.rf_ram.memory\[39\]\[7\] _01544_ _01545_ _02189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_91_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06591_ _02913_ _02914_ _02915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_75_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08330_ _03955_ _03956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_36_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05542_ _01492_ _02092_ _02101_ _02120_ _02121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_33_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09473__A2 _04711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08261_ _03703_ _03885_ _03891_ _00951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05473_ _01490_ _02043_ _02052_ _02053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__06287__A2 _02731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04917__S0 _01497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07212_ u_cpu.rf_ram.memory\[142\]\[4\] _03267_ _03272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08192_ u_arbiter.i_wb_cpu_dbus_dat\[12\] _03835_ _03848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09225__A2 _04563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07143_ _03110_ _03227_ _03233_ _00490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08984__A1 _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07787__A2 _03593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07074_ u_cpu.rf_ram.memory\[57\]\[7\] _03187_ _03195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05342__S0 _01523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05798__A1 _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06025_ u_cpu.cpu.ctrl.o_ibus_adr\[18\] _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_82_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07539__A2 _03455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07976_ _03697_ _03710_ _03713_ _00844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09715_ _00109_ io_in[4] u_cpu.rf_ram.memory\[21\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08478__C _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06927_ u_cpu.rf_ram.memory\[29\]\[6\] _03100_ _03113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05970__A1 _02418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09704__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05970__B2 u_arbiter.i_wb_cpu_dbus_adr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05183__B _01480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09646_ u_cpu.rf_ram.memory\[100\]\[4\] _04812_ _04817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06858_ u_cpu.rf_ram.memory\[66\]\[2\] _03069_ _03072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07711__A2 _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05809_ _02272_ u_cpu.rf_ram_if.rdata1\[5\] _02378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09577_ _04634_ _04772_ _04778_ _01380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05722__A1 _02259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06789_ u_cpu.rf_ram.memory\[75\]\[4\] _03028_ _03033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08528_ _03923_ _03918_ _04127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09854__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09464__A2 _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06278__A2 _02719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07475__A1 _03318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08459_ _01454_ _03956_ _04067_ _00973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10831__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09216__A2 _04563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08714__S _04257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10421_ _00794_ io_in[4] u_cpu.rf_ram.memory\[90\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07227__A1 _03104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07778__A2 _03593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10352_ _00738_ io_in[4] u_cpu.rf_ram.memory\[124\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05333__S0 _01497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10981__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06450__A2 _02829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10283_ _00669_ io_in[4] u_cpu.rf_ram.memory\[131\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10211__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07950__A2 _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09152__A1 _04448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07702__A2 _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10361__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09455__A2 _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06269__A2 _02719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05540__C _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06208__I _02641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09207__A2 _04553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10619_ _00992_ io_in[4] u_cpu.cpu.immdec.imm19_12_20\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05492__A3 _02071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07769__A2 _03583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05324__S0 _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06441__A2 _02816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09727__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08579__B _04164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07830_ _03508_ _03616_ _03623_ _00787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05252__I0 u_cpu.rf_ram.memory\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07941__A2 _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07761_ _03494_ _03583_ _03584_ _00757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_04973_ _01480_ _01558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10704__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06099__B _02313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09500_ _04724_ _04723_ _04731_ _01350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06712_ _02885_ _02988_ _02990_ _00302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07692_ u_cpu.rf_ram.memory\[125\]\[2\] _03543_ _03546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09877__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08497__A3 u_arbiter.i_wb_cpu_dbus_we vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09431_ u_cpu.rf_ram.memory\[86\]\[7\] _04681_ _04689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06643_ _02891_ _02945_ _02950_ _00273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05704__A1 _02259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09362_ _04650_ _04651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10854__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06574_ u_cpu.rf_ram.memory\[4\]\[3\] _02900_ _02904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_75_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09446__A2 _04691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08313_ u_arbiter.i_wb_cpu_rdt\[5\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[5\]
+ _02465_ _03941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07457__A1 _03318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05525_ u_cpu.rf_ram.memory\[32\]\[6\] u_cpu.rf_ram.memory\[33\]\[6\] u_cpu.rf_ram.memory\[34\]\[6\]
+ u_cpu.rf_ram.memory\[35\]\[6\] _01495_ _01499_ _02104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09293_ u_cpu.rf_ram.memory\[108\]\[5\] _04603_ _04609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08244_ u_arbiter.i_wb_cpu_rdt\[30\] _02924_ _03882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05456_ _01512_ _02035_ _02036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05022__I _01518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07209__A1 _03104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06680__A2 _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08175_ u_arbiter.i_wb_cpu_rdt\[6\] _03822_ _03833_ u_arbiter.i_wb_cpu_dbus_dat\[7\]
+ _03837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05387_ _01464_ _01967_ _01968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08957__A1 _03956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04861__I u_cpu.cpu.decode.op21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07126_ u_cpu.rf_ram.memory\[54\]\[6\] _03217_ _03224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05178__B _01558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06432__A2 _02816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07057_ _03114_ _03177_ _03185_ _00452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10234__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05893__S _02431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06008_ _02456_ _02513_ _02514_ _00074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_82_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09382__A1 _04622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06196__A1 _01460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07932__A2 _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10384__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07959_ _03701_ _03693_ _03702_ _00838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09134__A1 _04448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10970_ _01339_ io_in[4] u_cpu.rf_ram.memory\[87\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09685__A2 _04832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09629_ _04632_ _04802_ _04807_ _01403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06499__A2 _02851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09437__A2 _04691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07448__A1 u_cpu.rf_ram.memory\[49\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08645__B1 _04009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08496__I0 u_arbiter.i_wb_cpu_rdt\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07999__A2 _03720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06120__A1 _01460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05554__S0 _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08948__A1 _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10404_ _00777_ io_in[4] u_cpu.cpu.state.o_cnt_r\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10335_ _00721_ io_in[4] u_cpu.rf_ram.memory\[126\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06423__A2 _02805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10266_ _00652_ io_in[4] u_cpu.rf_ram.memory\[134\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10727__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10197_ _00583_ io_in[4] u_cpu.rf_ram.memory\[143\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07923__A2 _03672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10877__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09676__A2 _04832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__04946__I _01498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09428__A2 _04681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10107__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07439__A1 _03318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08100__A2 _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05310_ _01617_ _01891_ _01519_ _01892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06290_ _02632_ _02733_ _02734_ _00136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05545__S0 _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05241_ u_cpu.rf_ram.memory\[28\]\[3\] u_cpu.rf_ram.memory\[29\]\[3\] u_cpu.rf_ram.memory\[30\]\[3\]
+ u_cpu.rf_ram.memory\[31\]\[3\] _01497_ _01501_ _01823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06662__A2 _02956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10257__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08939__A1 _03932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08939__B2 _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05172_ _01543_ _01754_ _01755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09600__A2 _02754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06414__A2 _02805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09980_ _00374_ io_in[4] u_cpu.rf_ram.memory\[65\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08931_ _03932_ _03975_ _03988_ _03944_ _04188_ _04394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_115_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09364__A1 _02632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08167__A2 _03822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08862_ u_cpu.rf_ram.memory\[109\]\[3\] _04351_ _04355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06178__A1 u_cpu.rf_ram.memory\[82\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07813_ _02396_ u_cpu.cpu.state.o_cnt_r\[2\] _03614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__07914__A2 _03672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08793_ _04316_ _01058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_84_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09116__A1 _04448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07744_ u_cpu.rf_ram.memory\[38\]\[1\] _03573_ _03575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_04956_ _01540_ _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09667__A2 _04822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05017__I _01504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07675_ _03500_ _03533_ _03536_ _00719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04887_ u_cpu.cpu.immdec.imm19_12_20\[5\] u_cpu.rf_ram_if.rtrig0 _01474_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_80_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09414_ _04638_ _04671_ _04679_ _01316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06626_ u_cpu.rf_ram.memory\[16\]\[5\] _02935_ _02941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09419__A2 _04681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11032__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09345_ u_cpu.rf_ram.memory\[59\]\[0\] _04641_ _04642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06557_ _02656_ _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__04900__A2 _01438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05888__S _02418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05508_ _01506_ _02086_ _01481_ _02087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09276_ _04446_ _04593_ _04599_ _01258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06488_ _02669_ _02851_ _02852_ _00216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05536__S0 _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08642__A3 _04228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08227_ _03870_ _03871_ _00937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07850__A1 _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06653__A2 _02956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05439_ u_cpu.rf_ram.memory\[40\]\[5\] u_cpu.rf_ram.memory\[41\]\[5\] u_cpu.rf_ram.memory\[42\]\[5\]
+ u_cpu.rf_ram.memory\[43\]\[5\] _01551_ _01524_ _02019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_14_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05700__I1 _02276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08158_ u_arbiter.i_wb_cpu_dbus_dat\[4\] _02915_ _03823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_107_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07109_ _03112_ _03207_ _03214_ _00475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06405__A2 _02794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08089_ u_cpu.rf_ram.memory\[115\]\[5\] _03770_ _03776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09095__S _04485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10120_ _00514_ io_in[4] u_cpu.rf_ram.memory\[15\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08158__A2 _02915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10051_ _00445_ io_in[4] u_cpu.rf_ram.memory\[58\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06169__A1 _02611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07905__A2 _03662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05355__C _01560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09658__A2 _04822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10953_ _01322_ io_in[4] u_cpu.rf_ram.memory\[86\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10884_ _01253_ io_in[4] u_cpu.rf_ram.memory\[83\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06341__A1 _02691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06892__A2 _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08094__A1 _03707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05527__S0 _01551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06644__A2 _02945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08397__A2 _03904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10318_ _00704_ io_in[4] u_cpu.rf_ram.memory\[128\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09346__A1 _04622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05546__B _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10249_ _00635_ io_in[4] u_cpu.rf_ram.memory\[136\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05790_ _01445_ _02265_ _02364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09649__A2 _04812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11055__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08321__A2 _03948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07460_ u_cpu.rf_ram.memory\[49\]\[7\] _03405_ _03413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06411_ u_cpu.rf_ram.memory\[45\]\[1\] _02805_ _02807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06883__A2 _03079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07391_ _03374_ _03375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09915__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08592__B _04165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09130_ _04444_ _04513_ _04518_ _01193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06342_ u_cpu.rf_ram.memory\[80\]\[7\] _02756_ _02764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05518__S0 _01497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09061_ _04444_ _04476_ _04481_ _01161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06273_ u_cpu.rf_ram.memory\[20\]\[3\] _02719_ _02723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07832__A1 _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06635__A2 _02945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08012_ _02642_ _03730_ _03733_ _00860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05224_ _01621_ _01806_ _01807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09585__A1 _04622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08388__A2 _03956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05155_ u_cpu.rf_ram.memory\[24\]\[2\] u_cpu.rf_ram.memory\[25\]\[2\] u_cpu.rf_ram.memory\[26\]\[2\]
+ u_cpu.rf_ram.memory\[27\]\[2\] _01508_ _01509_ _01738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_144_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06399__A1 _02687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09963_ _00357_ io_in[4] u_cpu.rf_ram.memory\[67\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07060__A2 _03187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05086_ _01548_ _01669_ _01518_ _01670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_103_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08914_ u_cpu.rf_ram.memory\[93\]\[2\] _04381_ _04384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09894_ _00288_ io_in[4] u_cpu.rf_ram.memory\[119\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08845_ _04343_ _01083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08560__A2 _03908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08776_ u_cpu.rf_ram.memory\[30\]\[6\] _04299_ _04306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06571__A1 _02637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05988_ _02492_ _02486_ _02487_ _02498_ _02499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_26_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07727_ _03498_ _03563_ _03565_ _00742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_04939_ _01499_ _01524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10422__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07658_ u_cpu.rf_ram.memory\[127\]\[3\] _03523_ _03527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06609_ _01634_ _02929_ _02931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__06874__A2 _03079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07589_ _03484_ _03485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__04885__A1 _01466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09328_ _02646_ _04630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08076__A1 _03707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05509__S0 _01530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10572__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09259_ u_cpu.rf_ram.memory\[107\]\[6\] _04583_ _04590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06626__A2 _02935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08722__S _02335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08379__A2 _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11152_ _00086_ io_in[0] u_scanchain_local.module_data_in\[64\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07051__A2 _03177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10103_ _00497_ io_in[4] u_cpu.rf_ram.memory\[52\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05366__B _01946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11083_ u_cpu.rf_ram_if.wdata1_r\[7\] io_in[4] u_cpu.rf_ram_if.wdata1_r\[6\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08536__C1 _04131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08000__A1 _03703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10034_ _00428_ io_in[4] u_cpu.rf_ram.memory\[60\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11078__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06011__B1 _02398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08551__A2 _04052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06562__A1 _02895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05365__A2 _01936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09938__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10936_ _01305_ io_in[4] u_cpu.rf_ram.memory\[85\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05117__A2 _01700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06314__A1 _02642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10915__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10867_ _01236_ io_in[4] u_cpu.rf_ram.memory\[105\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05668__A3 _02245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06865__A2 _03069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04876__A1 _01439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10798_ _01167_ io_in[4] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06617__A2 _02935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07290__A2 _03308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09567__A1 _04622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05428__I0 u_cpu.rf_ram.memory\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07042__A2 _03177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08790__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06960_ u_cpu.rf_ram.memory\[62\]\[4\] _03127_ _03132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05911_ u_arbiter.i_wb_cpu_rdt\[26\] u_arbiter.i_wb_cpu_dbus_dat\[23\] _02431_ _02442_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_79_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06891_ _02881_ _03089_ _03090_ _00381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08587__B _03915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08630_ u_cpu.cpu.immdec.imm19_12_20\[8\] _03955_ _04219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10445__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05842_ _02388_ _02401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_27_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06553__A1 _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08561_ _04156_ _04157_ _04158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05773_ u_cpu.cpu.alu.i_rs1 u_cpu.cpu.alu.add_cy_r _02278_ _02348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_07512_ u_cpu.rf_ram.memory\[134\]\[6\] _03435_ _03442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05108__A2 _01691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08492_ _04000_ _04024_ _04055_ _04033_ _04095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_50_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10595__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07443_ _03322_ _03395_ _03403_ _00620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06856__A2 _03069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05903__I1 u_arbiter.i_wb_cpu_dbus_dat\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08058__A1 _03707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07374_ u_cpu.rf_ram.memory\[14\]\[0\] _03365_ _03366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09113_ u_cpu.rf_ram.memory\[101\]\[5\] _04503_ _04509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06069__B1 _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06325_ _02614_ _02716_ _02754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06608__A2 _02929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09044_ _04450_ _04463_ _04471_ _01154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06256_ _02687_ _02707_ _02712_ _00124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06126__I _02606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07281__A2 _03308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05207_ _01554_ _01789_ _01607_ _01790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_117_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06187_ _02664_ _02368_ _02611_ _02665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05138_ _01512_ _01721_ _01481_ _01722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07033__A2 _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05069_ u_cpu.rf_ram.memory\[20\]\[1\] u_cpu.rf_ram.memory\[21\]\[1\] u_cpu.rf_ram.memory\[22\]\[1\]
+ u_cpu.rf_ram.memory\[23\]\[1\] _01497_ _01501_ _01653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09946_ _00340_ io_in[4] u_cpu.rf_ram.memory\[75\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06792__A1 _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09877_ _00271_ io_in[4] u_cpu.rf_ram.memory\[17\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08533__A2 _04131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08828_ u_cpu.cpu.ctrl.o_ibus_adr\[21\] _04327_ _04329_ u_cpu.cpu.ctrl.o_ibus_adr\[22\]
+ _04335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_100_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06544__A1 _02881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08759_ _04288_ _04295_ _04296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10938__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10721_ _01091_ io_in[4] u_cpu.rf_ram.memory\[109\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06847__A2 _03059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10652_ _01025_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09097__I0 u_arbiter.i_wb_cpu_rdt\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04953__S1 _01532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10583_ _00956_ io_in[4] u_cpu.cpu.decode.opcode\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08960__B _03948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07272__A2 _03297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10318__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09549__A1 _04622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07024__A2 _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08772__A2 _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11135_ _00067_ io_in[0] u_scanchain_local.module_data_in\[47\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10468__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11066_ u_cpu.rf_ram_if.wdata0_r\[3\] io_in[4] u_cpu.rf_ram_if.wdata0_r\[2\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09760__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08524__A2 _04101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10017_ _00411_ io_in[4] u_cpu.rf_ram.memory\[62\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06535__A1 _02689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08288__A1 _02465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06838__A2 _03059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10919_ _01288_ io_in[4] u_cpu.rf_ram.memory\[59\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05197__S1 _01531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05897__I0 u_arbiter.i_wb_cpu_rdt\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06110_ _02259_ _02598_ _02599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07263__A2 _03297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08460__A1 _02265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07090_ u_cpu.rf_ram.memory\[56\]\[6\] _03197_ _03204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06041_ _02456_ _02541_ _02542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07015__A2 _03157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09800_ _00194_ io_in[4] u_cpu.rf_ram.memory\[44\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07992_ _03695_ _03720_ _03722_ _00851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06774__A1 _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09731_ _00125_ io_in[4] u_cpu.rf_ram.memory\[18\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06943_ _03108_ _03117_ _03122_ _00401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09662_ u_cpu.rf_ram.memory\[89\]\[3\] _04822_ _04826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06874_ u_cpu.rf_ram.memory\[65\]\[1\] _03079_ _03081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08613_ _04013_ _04052_ _04179_ _04203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05825_ _01467_ _02377_ _02386_ _00013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09593_ _04632_ _04782_ _04787_ _01387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_43_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08544_ u_cpu.cpu.immdec.imm30_25\[5\] _04104_ _04142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08279__A1 _02465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05756_ _02330_ _02331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08475_ _03906_ _04079_ _04080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06829__A2 _03049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05687_ u_cpu.cpu.immdec.imm11_7\[0\] _02264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_51_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05888__I0 u_arbiter.i_wb_cpu_rdt\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07426_ _02838_ _02976_ _03394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09079__I0 u_arbiter.i_wb_cpu_rdt\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05501__A2 _02080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07357_ _03306_ _03355_ _03356_ _00581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08780__B _02395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06308_ _02744_ _02745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08272__S _02465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08451__A1 _03925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07254__A2 _03287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07288_ _02651_ _03316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08451__B2 _03941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09027_ _02754_ _04349_ _04462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06239_ u_cpu.rf_ram.memory\[81\]\[5\] _02697_ _02703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05360__S1 _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10610__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07006__A2 _03157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05628__C _01485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09783__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08754__A2 u_cpu.cpu.state.o_cnt_r\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05112__S1 _01594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09929_ _00323_ io_in[4] u_cpu.rf_ram.memory\[74\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10760__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11084__D u_cpu.cpu.o_wdata1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08955__B _03923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11116__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05740__A2 u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10704_ _01074_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07493__A2 _03425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10140__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10635_ _01008_ io_in[4] u_cpu.rf_ram.memory\[31\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08442__A1 _03906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10566_ _00939_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07245__A2 _03287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08993__A2 _04436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10497_ _00870_ io_in[4] u_cpu.rf_ram.memory\[11\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10290__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05351__S1 _01524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05103__S1 _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05559__A2 _02137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06756__A1 _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11118_ _00049_ io_in[0] u_arbiter.i_wb_cpu_rdt\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11049_ _01418_ io_in[4] u_cpu.rf_ram.memory\[89\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04949__I _01519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06508__A1 _02681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09170__A2 _04533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07181__A1 _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05610_ _02181_ _02183_ _02185_ _02187_ _01541_ _02188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_64_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06590_ _02307_ _02311_ _02914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05541_ _01490_ _02110_ _02119_ _02120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_08260_ u_cpu.rf_ram.memory\[113\]\[5\] _03885_ _03891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05472_ _02045_ _02047_ _02049_ _02051_ _01581_ _02052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__07484__A2 _03425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04917__S1 _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07211_ _03106_ _03267_ _03271_ _00520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05495__A1 _01465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08191_ _03846_ _03847_ _00925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10633__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07142_ u_cpu.rf_ram.memory\[53\]\[5\] _03227_ _03233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07236__A2 _03277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05098__I1 u_cpu.rf_ram.memory\[49\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08984__A2 _02766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07073_ _03112_ _03187_ _03194_ _00459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05798__A2 _02369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06995__A1 _03106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05342__S1 _01525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06024_ _02463_ _02526_ _02527_ _00077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10783__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07975_ u_cpu.rf_ram.memory\[118\]\[2\] _03710_ _03713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09714_ _00108_ io_in[4] u_cpu.rf_ram.memory\[21\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10013__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06926_ _02661_ _03112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11139__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09161__A2 _04533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09645_ _04630_ _04812_ _04816_ _01410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06857_ _02885_ _03069_ _03071_ _00366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05808_ _02273_ u_cpu.rf_ram.rdata\[5\] _02377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09576_ u_cpu.rf_ram.memory\[25\]\[5\] _04772_ _04778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06788_ _02889_ _03028_ _03032_ _00336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10163__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08527_ _04123_ _04126_ _00982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05739_ _02313_ _01441_ _02314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_23_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08458_ _04009_ _04050_ _04064_ _04066_ _04067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08672__A1 _03691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07475__A2 _03415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05486__A1 _01617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07409_ _03384_ _03385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05030__S0 _01496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08389_ _03895_ _03965_ _04009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10420_ _00793_ io_in[4] u_cpu.rf_ram.memory\[90\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07227__A2 _03277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08975__A2 _04425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10351_ _00737_ io_in[4] u_cpu.rf_ram.memory\[124\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05333__S1 _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06986__A1 _02814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10282_ _00668_ io_in[4] u_cpu.rf_ram.memory\[132\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08730__S _02335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06738__A1 _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05374__B _01558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05961__A2 _02461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09152__A2 _04523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10506__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07163__A1 _03112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06910__A1 _03098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10656__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07466__A2 _03415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05477__A1 _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05021__S0 _01576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08415__A1 _03935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07218__A2 _03267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10618_ _00991_ io_in[4] u_cpu.cpu.immdec.imm19_12_20\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05229__A1 _01792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10549_ _00922_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05324__S1 _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06977__A1 _03106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10036__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09391__A2 _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07760_ u_cpu.rf_ram.memory\[37\]\[0\] _03583_ _03584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04972_ u_cpu.rf_ram.memory\[44\]\[0\] u_cpu.rf_ram.memory\[45\]\[0\] u_cpu.rf_ram.memory\[46\]\[0\]
+ u_cpu.rf_ram.memory\[47\]\[0\] _01555_ _01556_ _01557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_56_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09143__A2 _04523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06711_ u_cpu.rf_ram.memory\[139\]\[1\] _02988_ _02990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10186__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07691_ _03498_ _03543_ _03545_ _00726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09430_ _04636_ _04681_ _04688_ _01323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06642_ u_cpu.rf_ram.memory\[17\]\[4\] _02945_ _02950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06901__A1 _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09361_ _02731_ _02780_ _04650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06573_ _02642_ _02900_ _02903_ _00250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_40_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08312_ u_arbiter.i_wb_cpu_rdt\[6\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[6\]
+ _02465_ _03940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05524_ _01571_ _02102_ _02103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09292_ _04444_ _04603_ _04608_ _01265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08654__A1 _03691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07457__A2 _03405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08243_ _02450_ _03874_ _03881_ _00943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05455_ u_cpu.rf_ram.memory\[100\]\[5\] u_cpu.rf_ram.memory\[101\]\[5\] u_cpu.rf_ram.memory\[102\]\[5\]
+ u_cpu.rf_ram.memory\[103\]\[5\] _01551_ _01524_ _02035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_119_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08174_ u_arbiter.i_wb_cpu_dbus_dat\[6\] _03835_ _03836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08406__A1 _03974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07209__A2 _03267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05386_ u_cpu.rf_ram.memory\[92\]\[4\] u_cpu.rf_ram.memory\[93\]\[4\] u_cpu.rf_ram.memory\[94\]\[4\]
+ u_cpu.rf_ram.memory\[95\]\[4\] _01562_ _01563_ _01967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07125_ _03110_ _03217_ _03223_ _00482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08957__A2 _04417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06968__A1 _02803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07056_ u_cpu.rf_ram.memory\[58\]\[7\] _03177_ _03185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06007_ _02418_ u_scanchain_local.module_data_in\[52\] _02398_ u_arbiter.i_wb_cpu_dbus_adr\[15\]
+ _02514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_114_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09382__A2 _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10529__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07393__A1 _03306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05194__B _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07958_ u_cpu.rf_ram.memory\[120\]\[4\] _03693_ _03702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09821__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09134__A2 _04513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06909_ u_cpu.rf_ram.memory\[29\]\[0\] _03100_ _03101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07145__A1 _03112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07889_ _02782_ _02825_ _03661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09628_ u_cpu.rf_ram.memory\[98\]\[4\] _04802_ _04807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10679__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07696__A2 _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08893__A1 _02632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09559_ _04634_ _04762_ _04768_ _01372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_19_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09971__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08645__A1 u_cpu.cpu.immdec.imm31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07448__A2 _03405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08496__I1 u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05554__S1 _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10403_ _00776_ io_in[4] u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10059__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06959__A1 _03106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10334_ _00720_ io_in[4] u_cpu.rf_ram.memory\[126\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10265_ _00651_ io_in[4] u_cpu.rf_ram.memory\[134\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09373__A2 _04651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10196_ _00582_ io_in[4] u_cpu.rf_ram.memory\[143\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09125__A2 _04513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05551__C _01560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08636__A1 _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07439__A2 _03395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05545__S1 _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05240_ _01473_ _01773_ _01822_ _00002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08939__A2 _04009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05171_ u_cpu.rf_ram.memory\[36\]\[2\] u_cpu.rf_ram.memory\[37\]\[2\] u_cpu.rf_ram.memory\[38\]\[2\]
+ u_cpu.rf_ram.memory\[39\]\[2\] _01544_ _01545_ _01754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09061__A1 _04444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08930_ _03932_ _03939_ _03948_ _03962_ _04393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_112_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09844__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09364__A2 _04651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08861_ _03697_ _04351_ _04354_ _01088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07375__A1 _02632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06178__A2 _02628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07812_ _02395_ _02359_ _00779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08792_ u_cpu.cpu.ctrl.o_ibus_adr\[4\] _04309_ _04311_ u_cpu.cpu.ctrl.o_ibus_adr\[5\]
+ _04316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10821__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09116__A2 _04503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07743_ _03494_ _03573_ _03574_ _00749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_04955_ _01483_ _01484_ _01540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07127__A1 _03112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09994__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08324__B1 _03915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07674_ u_cpu.rf_ram.memory\[126\]\[2\] _03533_ _03536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07678__A2 _03533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04886_ _01472_ _01473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08875__A1 _02632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05689__A1 _01444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09413_ u_cpu.rf_ram.memory\[110\]\[7\] _04671_ _04679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06625_ _02891_ _02935_ _02940_ _00265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10971__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06350__A2 _02770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08627__A1 _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06556_ _02891_ _02883_ _02892_ _00244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09344_ _04640_ _04641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05507_ u_cpu.rf_ram.memory\[24\]\[6\] u_cpu.rf_ram.memory\[25\]\[6\] u_cpu.rf_ram.memory\[26\]\[6\]
+ u_cpu.rf_ram.memory\[27\]\[6\] _01522_ _01509_ _02086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_139_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09275_ u_cpu.rf_ram.memory\[83\]\[5\] _04593_ _04599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06487_ u_cpu.rf_ram.memory\[43\]\[0\] _02851_ _02852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10201__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05536__S1 _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08226_ u_arbiter.i_wb_cpu_rdt\[23\] _03807_ _03829_ u_arbiter.i_wb_cpu_dbus_dat\[24\]
+ _03871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_138_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05438_ _01504_ _02017_ _01518_ _02018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_101_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07850__A2 _03626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05861__A1 _02414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08157_ _03807_ _03822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05369_ u_cpu.rf_ram.memory\[96\]\[4\] u_cpu.rf_ram.memory\[97\]\[4\] u_cpu.rf_ram.memory\[98\]\[4\]
+ u_cpu.rf_ram.memory\[99\]\[4\] _01567_ _01568_ _01950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_101_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07108_ u_cpu.rf_ram.memory\[55\]\[6\] _03207_ _03214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08088_ _03701_ _03770_ _03775_ _00894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07602__A2 _03485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10351__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07039_ _02667_ _03167_ _03175_ _00444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_134_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10050_ _00444_ io_in[4] u_cpu.rf_ram.memory\[5\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09355__A2 _04641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09107__A2 _04503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10952_ _01321_ io_in[4] u_cpu.rf_ram.memory\[86\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10883_ _01252_ io_in[4] u_cpu.rf_ram.memory\[107\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06341__A2 _02756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09717__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08094__A2 _03770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05527__S1 _01524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07841__A2 _03626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05852__A1 _02355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05099__B _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09867__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09594__A2 _04782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10317_ _00703_ io_in[4] u_cpu.rf_ram.memory\[128\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10844__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09346__A2 _04641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10248_ _00634_ io_in[4] u_cpu.rf_ram.memory\[136\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07357__A1 _03306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10179_ _00565_ io_in[4] u_cpu.rf_ram.memory\[71\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10994__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07109__A1 _03112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06580__A2 _02900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08857__A1 _03691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06332__A2 _02756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06410_ _02669_ _02805_ _02806_ _00184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10224__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08609__A1 _04165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07390_ _02780_ _02976_ _03374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06341_ _02691_ _02756_ _02763_ _00158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08085__A2 _03770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05518__S1 _01525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06096__A1 u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09060_ u_cpu.rf_ram.memory\[28\]\[4\] _04476_ _04481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06272_ _02683_ _02719_ _02722_ _00130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07832__A2 _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10374__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08011_ u_cpu.rf_ram.memory\[8\]\[2\] _03730_ _03733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05223_ u_cpu.rf_ram.memory\[72\]\[2\] u_cpu.rf_ram.memory\[73\]\[2\] u_cpu.rf_ram.memory\[74\]\[2\]
+ u_cpu.rf_ram.memory\[75\]\[2\] _01522_ _01622_ _01806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09034__A1 _04440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09585__A2 _04782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05154_ _01493_ _01736_ _01737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06399__A2 _02794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05085_ u_cpu.rf_ram.memory\[32\]\[1\] u_cpu.rf_ram.memory\[33\]\[1\] u_cpu.rf_ram.memory\[34\]\[1\]
+ u_cpu.rf_ram.memory\[35\]\[1\] _01495_ _01499_ _01669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09962_ _00356_ io_in[4] u_cpu.rf_ram.memory\[68\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08913_ _03695_ _04381_ _04383_ _01111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09893_ _00287_ io_in[4] u_cpu.rf_ram.memory\[119\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08844_ u_cpu.cpu.ctrl.o_ibus_adr\[29\] _04327_ _04329_ u_cpu.cpu.ctrl.o_ibus_adr\[30\]
+ _04343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_44_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07899__A2 _03662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06020__A1 _02389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08775_ _03703_ _04299_ _04305_ _01051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05987_ u_cpu.cpu.ctrl.o_ibus_adr\[11\] u_cpu.cpu.ctrl.o_ibus_adr\[10\] _02498_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06571__A2 _02900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07726_ u_cpu.rf_ram.memory\[123\]\[1\] _03563_ _03565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04938_ _01522_ _01523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__04867__I u_cpu.cpu.decode.op26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05206__S0 _01576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07657_ _03500_ _03523_ _03526_ _00711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_04869_ _01447_ _01449_ _01456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_13_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06323__A2 _02745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05899__S _02431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06608_ _01634_ _02929_ _02930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07588_ _02731_ _02814_ _03484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09327_ _04628_ _04624_ _04629_ _01279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10717__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04885__A2 _01471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06539_ _02693_ _02872_ _02880_ _00239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08076__A2 _03760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05509__S1 _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09258_ _04446_ _04583_ _04589_ _01250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07823__A2 _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05834__A1 _01444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08209_ _03858_ _03859_ _00931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09189_ u_cpu.rf_ram.memory\[99\]\[7\] _04543_ _04551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10867__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09576__A2 _04772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07587__A1 _03322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08784__B1 _04311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11151_ _00085_ io_in[0] u_scanchain_local.module_data_in\[63\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05647__B _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10102_ _00496_ io_in[4] u_cpu.rf_ram.memory\[52\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11082_ u_cpu.rf_ram_if.wdata1_r\[6\] io_in[4] u_cpu.rf_ram_if.wdata1_r\[5\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07339__A1 _03306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08536__C2 _03959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10033_ _00427_ io_in[4] u_cpu.rf_ram.memory\[60\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07862__B _01441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08000__A2 _03720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06011__A1 _02418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06562__A2 _02883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05365__A3 _01945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10247__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09500__A2 _04723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10935_ _01304_ io_in[4] u_cpu.rf_ram.memory\[85\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06314__A2 _02745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07511__A1 _03318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10866_ _01235_ io_in[4] u_cpu.rf_ram.memory\[105\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10397__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04876__A2 _01438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08067__A2 _03760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10797_ _01166_ io_in[4] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06078__A1 _02456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05825__A1 _01467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09016__A1 _04440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09567__A2 _04772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06250__A1 _02681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05276__C _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11022__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08378__I0 u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05910_ _02441_ _00046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06890_ u_cpu.rf_ram.memory\[64\]\[0\] _03089_ _03090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06002__A1 u_cpu.cpu.ctrl.o_ibus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05841_ u_arbiter.i_wb_cpu_dbus_we _02400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_94_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06553__A2 _02883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08560_ _03899_ _03908_ _03909_ _03925_ _04031_ _04157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_05772_ u_cpu.cpu.bne_or_bge _02344_ _02345_ _02346_ _02347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_48_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07511_ _03318_ _03435_ _03441_ _00650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_63_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08491_ _03963_ _04093_ _03899_ _04094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07442_ u_cpu.rf_ram.memory\[137\]\[7\] _03395_ _03403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05513__B1 _02089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07373_ _03364_ _03365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08058__A2 _03750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06069__A1 _02402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09112_ _04444_ _04503_ _04508_ _01185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06324_ _02667_ _02745_ _02753_ _00151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_108_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09043_ u_cpu.rf_ram.memory\[96\]\[7\] _04463_ _04471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06255_ u_cpu.rf_ram.memory\[18\]\[4\] _02707_ _02712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05206_ u_cpu.rf_ram.memory\[116\]\[2\] u_cpu.rf_ram.memory\[117\]\[2\] u_cpu.rf_ram.memory\[118\]\[2\]
+ u_cpu.rf_ram.memory\[119\]\[2\] _01576_ _01577_ _01789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09558__A2 _04762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06186_ u_cpu.rf_ram_if.wdata1_r\[7\] _02664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_132_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07569__A1 _03322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05137_ u_cpu.rf_ram.memory\[76\]\[1\] u_cpu.rf_ram.memory\[77\]\[1\] u_cpu.rf_ram.memory\[78\]\[1\]
+ u_cpu.rf_ram.memory\[79\]\[1\] _01529_ _01500_ _01721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__05467__B _01600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05068_ _01506_ _01651_ _01481_ _01652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09945_ _00339_ io_in[4] u_cpu.rf_ram.memory\[75\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08518__B1 _03988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06792__A2 _03028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09876_ _00270_ io_in[4] u_cpu.rf_ram.memory\[17\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08827_ _04334_ _01074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06544__A2 _02883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08758_ u_arbiter.i_wb_cpu_dbus_adr\[2\] _02598_ _04295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07709_ _03498_ _03553_ _03555_ _00734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_54_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08689_ _02335_ _04257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09494__A1 u_cpu.cpu.state.genblk1.misalign_trap_sync_r vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10720_ _01090_ io_in[4] u_cpu.rf_ram.memory\[109\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08049__A2 _03750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10651_ _01024_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10582_ _00955_ io_in[4] u_cpu.cpu.decode.opcode\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08960__C _04031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05807__A1 _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09549__A2 _04762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11045__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05035__A2 _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06232__A1 _02681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11134_ _00066_ io_in[0] u_scanchain_local.module_data_in\[46\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07980__A1 _03701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06783__A2 _03028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09905__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11065_ u_cpu.rf_ram_if.wdata0_r\[2\] io_in[4] u_cpu.rf_ram_if.wdata0_r\[1\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05991__B1 _02398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10016_ _00410_ io_in[4] u_cpu.rf_ram.memory\[62\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06535__A2 _02872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08532__I0 u_arbiter.i_wb_cpu_rdt\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10918_ _01287_ io_in[4] u_cpu.rf_ram.memory\[59\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07611__I _02636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05897__I1 u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10849_ _01218_ io_in[4] u_cpu.rf_ram.memory\[99\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08643__S _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07799__A1 _02395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08460__A2 _02400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06040_ u_cpu.cpu.ctrl.o_ibus_adr\[21\] _02539_ _02541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06471__A1 _02681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04970__I _01494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10412__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07991_ u_cpu.rf_ram.memory\[121\]\[1\] _03720_ _03722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06774__A2 _03018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08598__B _03975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09730_ _00124_ io_in[4] u_cpu.rf_ram.memory\[18\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06942_ u_cpu.rf_ram.memory\[63\]\[4\] _03117_ _03122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05982__B1 _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09661_ _04628_ _04822_ _04825_ _01417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06873_ _02881_ _03079_ _03080_ _00373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10562__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06526__A2 _02872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08612_ _02909_ _02411_ _04201_ _04202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05824_ u_cpu.rf_ram_if.rdata0\[6\] _01467_ _02386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09592_ u_cpu.rf_ram.memory\[24\]\[4\] _04782_ _04787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08543_ _04009_ _04136_ _04140_ _03955_ _04141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05755_ _02266_ _02326_ _02329_ u_arbiter.i_wb_cpu_ibus_adr\[0\] _02330_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__09476__A1 _04628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08279__A2 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08474_ _03996_ _03908_ _04079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05686_ u_cpu.cpu.bufreg2.i_cnt_done _02263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_126_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07425_ _03322_ _03385_ _03393_ _00612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07356_ u_cpu.rf_ram.memory\[143\]\[0\] _03355_ _03356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11068__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06307_ _02731_ _02743_ _02744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07287_ _03314_ _03308_ _03315_ _00552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08451__A2 _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09026_ _04450_ _04453_ _04461_ _01146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__04880__I _01438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06462__A1 _02691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06238_ _02687_ _02697_ _02702_ _00116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08352__I _03963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09928__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06169_ _02611_ u_cpu.rf_ram_if.wdata0_r\[4\] _02649_ _02650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10092__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09400__A1 _04622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07962__A1 _03703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06765__A2 _03018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10905__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09928_ _00322_ io_in[4] u_cpu.rf_ram.memory\[74\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09859_ _00253_ io_in[4] u_cpu.rf_ram.memory\[4\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06517__A2 _02861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08728__S _02335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07190__A2 _03257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10703_ _01073_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10634_ _01007_ io_in[4] u_cpu.rf_ram.memory\[31\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08442__A2 _03947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10565_ _00938_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10435__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10496_ _00869_ io_in[4] u_cpu.rf_ram.memory\[11\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05008__A2 _01588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10585__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07953__A1 _03697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06756__A2 _03008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11117_ _00047_ io_in[0] u_arbiter.i_wb_cpu_rdt\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07606__I _02631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11048_ _01417_ io_in[4] u_cpu.rf_ram.memory\[89\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06508__A2 _02861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07181__A2 _03247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05192__A1 _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09458__A1 _04628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05540_ _02112_ _02114_ _02116_ _02118_ _01581_ _02119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_51_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08130__A1 _03707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05471_ _01554_ _02050_ _01607_ _02051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_60_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08681__A2 _04247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07210_ u_cpu.rf_ram.memory\[142\]\[3\] _03267_ _03271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08190_ u_arbiter.i_wb_cpu_rdt\[11\] _03822_ _03833_ u_arbiter.i_wb_cpu_dbus_dat\[12\]
+ _03847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__05495__A2 _02074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06692__A1 _02881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07141_ _03108_ _03227_ _03232_ _00489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08433__A2 _04041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07072_ u_cpu.rf_ram.memory\[57\]\[6\] _03187_ _03194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06023_ _02402_ u_scanchain_local.module_data_in\[55\] _02478_ u_arbiter.i_wb_cpu_dbus_adr\[18\]
+ _02527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10928__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06995__A2 _03147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07944__A1 _02954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06747__A2 _03008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07974_ _03695_ _03710_ _03712_ _00843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09713_ _00107_ io_in[4] u_cpu.rf_ram.memory\[21\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06925_ _03110_ _03100_ _03111_ _00394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09697__A1 _02396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09644_ u_cpu.rf_ram.memory\[100\]\[3\] _04812_ _04816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06856_ u_cpu.rf_ram.memory\[66\]\[1\] _03069_ _03071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05036__I _01504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07172__A2 _03247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10308__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05807_ _02272_ _02375_ _02376_ _00018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_82_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09575_ _04632_ _04772_ _04777_ _01379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05183__A1 _01566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06787_ u_cpu.rf_ram.memory\[75\]\[3\] _03028_ _03032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08526_ u_cpu.cpu.immdec.imm30_25\[3\] _04102_ _04124_ u_cpu.cpu.immdec.imm30_25\[4\]
+ _04125_ _03959_ _04126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XANTENNA__04930__A1 _01513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05738_ _01444_ _02313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_35_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08457_ _03910_ _04065_ _03966_ _04066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05669_ _02227_ _02246_ _01471_ _02247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08672__A2 _04247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10458__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06683__A1 _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05486__A2 _02065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07408_ _02743_ _02782_ _03384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05030__S1 _01594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08388_ _02309_ _03956_ _04008_ _00961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05700__S u_arbiter.i_wb_cpu_dbus_we vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07339_ _03306_ _03345_ _03346_ _00573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09750__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09621__A1 _04622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06435__A1 _02685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10350_ _00736_ io_in[4] u_cpu.rf_ram.memory\[124\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05639__C _01560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06986__A2 _02827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09009_ _02626_ _02870_ _04452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10281_ _00667_ io_in[4] u_cpu.rf_ram.memory\[132\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06738__A2 _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08360__A1 _03950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07163__A2 _03237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05174__A1 _01548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06910__A2 _03100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08112__A1 _03707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08663__A2 _04237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05021__S1 _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10617_ _00990_ io_in[4] u_cpu.cpu.csr_imm vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09612__A1 u_cpu.rf_ram.memory\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06426__A1 _02782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10548_ _00921_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06977__A2 _03137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10479_ _00852_ io_in[4] u_cpu.rf_ram.memory\[121\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06729__A2 _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05565__B _01600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09679__A1 _04628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04971_ _01498_ _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_49_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06710_ _02881_ _02988_ _02989_ _00301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_77_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07690_ u_cpu.rf_ram.memory\[125\]\[1\] _03543_ _03545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07154__A2 _03237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06641_ _02889_ _02945_ _02949_ _00272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05165__A1 _01528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06901__A2 _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09360_ _04638_ _04641_ _04649_ _01292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06572_ u_cpu.rf_ram.memory\[4\]\[2\] _02900_ _02903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10600__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08311_ _03901_ _03938_ _03939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_75_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05523_ u_cpu.rf_ram.memory\[36\]\[6\] u_cpu.rf_ram.memory\[37\]\[6\] u_cpu.rf_ram.memory\[38\]\[6\]
+ u_cpu.rf_ram.memory\[39\]\[6\] _01544_ _01545_ _02102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09291_ u_cpu.rf_ram.memory\[108\]\[4\] _04603_ _04608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09773__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08654__A2 _04237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08242_ u_arbiter.i_wb_cpu_rdt\[29\] _03807_ _03808_ u_arbiter.i_wb_cpu_dbus_dat\[29\]
+ _03881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05454_ _01492_ _02005_ _02014_ _02033_ _02034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_123_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10750__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05385_ _01490_ _01956_ _01965_ _01966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_08173_ _03808_ _03835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08406__A2 _04024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09603__A1 _02669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07124_ u_cpu.rf_ram.memory\[54\]\[5\] _03217_ _03223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06968__A2 _02827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07055_ _03112_ _03177_ _03184_ _00451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11106__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06006_ u_cpu.cpu.ctrl.o_ibus_adr\[15\] _02512_ _02513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_47_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08590__A1 _03965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07393__A2 _03375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06196__A3 _02612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10130__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07957_ _02651_ _03701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_75_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06908_ _03099_ _03100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07888_ _03510_ _03652_ _03660_ _00809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07145__A2 _03227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09627_ _04630_ _04802_ _04806_ _01402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_16_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05156__A1 _01506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06839_ _02885_ _03059_ _03061_ _00358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_16_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08893__A2 _04371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10280__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09558_ u_cpu.rf_ram.memory\[26\]\[5\] _04762_ _04768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08509_ _03901_ _04095_ _04108_ _04109_ _04110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__08645__A2 _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09489_ _04720_ _04721_ _04722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_11_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06656__A1 _02885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10402_ _00775_ io_in[4] u_cpu.cpu.mem_bytecnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06959__A2 _03127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07081__A1 _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10333_ _00719_ io_in[4] u_cpu.rf_ram.memory\[126\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10264_ _00650_ io_in[4] u_cpu.rf_ram.memory\[134\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10195_ _00581_ io_in[4] u_cpu.rf_ram.memory\[143\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08581__A1 _04000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07384__A2 _03365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10623__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08333__A1 _02911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04993__I1 u_cpu.rf_ram.memory\[49\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07136__A2 _03227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05147__A1 _01465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09796__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08884__A2 _04361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06895__A1 _02887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05698__A2 _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10773__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08636__A2 u_arbiter.i_wb_cpu_rdt\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06647__A1 _02895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10003__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11129__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05170_ _01746_ _01748_ _01750_ _01752_ _01541_ _01753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__09061__A2 _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10153__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05295__B _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08860_ u_cpu.rf_ram.memory\[109\]\[2\] _04351_ _04354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07375__A2 _03365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07811_ _03613_ _00778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_111_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08791_ _04315_ _01057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_07742_ u_cpu.rf_ram.memory\[38\]\[0\] _03573_ _03574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04954_ _01513_ _01538_ _01482_ _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_42_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08324__A1 _03899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07127__A2 _03217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05138__A1 _01512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07673_ _03498_ _03533_ _03535_ _00718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_04885_ _01466_ _01471_ _01472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08875__A2 _04361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09412_ _04636_ _04671_ _04678_ _01315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06624_ u_cpu.rf_ram.memory\[16\]\[4\] _02935_ _02940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05689__A2 _02265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09343_ _02827_ _02849_ _04640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06555_ u_cpu.rf_ram.memory\[50\]\[4\] _02883_ _02892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08627__A2 u_arbiter.i_wb_cpu_rdt\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05506_ _01493_ _02084_ _02085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09274_ _04444_ _04593_ _04598_ _01257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06486_ _02850_ _02851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08225_ u_arbiter.i_wb_cpu_dbus_dat\[23\] _03808_ _03870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05310__A1 _01617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05437_ u_cpu.rf_ram.memory\[32\]\[5\] u_cpu.rf_ram.memory\[33\]\[5\] u_cpu.rf_ram.memory\[34\]\[5\]
+ u_cpu.rf_ram.memory\[35\]\[5\] _01495_ _01499_ _02017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_20_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05368_ _01571_ _01948_ _01949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05861__A2 _02403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08156_ _03821_ _00916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_140_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09052__A2 _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07107_ _03110_ _03207_ _03213_ _00474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07063__A1 _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08087_ u_cpu.rf_ram.memory\[115\]\[4\] _03770_ _03775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05299_ _01464_ _01880_ _01881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07038_ u_cpu.rf_ram.memory\[5\]\[7\] _03167_ _03175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_88_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10646__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08563__A1 _03925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07366__A2 _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05377__A1 _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08989_ u_cpu.rf_ram.memory\[94\]\[1\] _04436_ _04439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08315__A1 _02465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07118__A2 _03217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10951_ _01320_ io_in[4] u_cpu.rf_ram.memory\[86\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05129__A1 _01617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10796__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08866__A2 _04351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06877__A1 _02887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10882_ _01251_ io_in[4] u_cpu.rf_ram.memory\[107\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08736__S _02335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10026__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06629__A1 _02895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09291__A2 _04603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05301__A1 _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10176__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09043__A2 _04463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06801__A1 _02632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10316_ _00702_ io_in[4] u_cpu.rf_ram.memory\[128\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10247_ _00633_ io_in[4] u_cpu.rf_ram.memory\[136\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08554__A1 _03925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07357__A2 _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08554__B2 _03908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05368__A1 _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10178_ _00564_ io_in[4] u_cpu.rf_ram.memory\[73\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08306__A1 _02466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07109__A2 _03207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07614__I _02641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08857__A2 _04351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05915__I0 u_arbiter.i_wb_cpu_rdt\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08609__A2 _04197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04973__I _01480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06340_ u_cpu.rf_ram.memory\[80\]\[6\] _02756_ _02763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10519__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06271_ u_cpu.rf_ram.memory\[20\]\[2\] _02719_ _02722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07293__A1 _03318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05222_ _01617_ _01804_ _01519_ _01805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08010_ _02637_ _03730_ _03732_ _00859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09811__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09034__A2 _04463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05153_ u_cpu.rf_ram.memory\[28\]\[2\] u_cpu.rf_ram.memory\[29\]\[2\] u_cpu.rf_ram.memory\[30\]\[2\]
+ u_cpu.rf_ram.memory\[31\]\[2\] _01497_ _01501_ _01736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07045__A1 _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08242__B1 _03808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10669__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07596__A2 _03485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05084_ _01543_ _01667_ _01668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09961_ _00355_ io_in[4] u_cpu.rf_ram.memory\[68\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08912_ u_cpu.rf_ram.memory\[93\]\[1\] _04381_ _04383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09961__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09892_ _00286_ io_in[4] u_cpu.rf_ram.memory\[119\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07348__A2 _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08843_ _04342_ _01082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05359__A1 _01566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08774_ u_cpu.rf_ram.memory\[30\]\[5\] _04299_ _04305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05986_ _02463_ _02496_ _02497_ _00068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07725_ _03494_ _03563_ _03564_ _00741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05472__C _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04937_ _01495_ _01522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_72_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10049__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06859__A1 _02887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05206__S1 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07656_ u_cpu.rf_ram.memory\[127\]\[2\] _03523_ _03526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04868_ u_cpu.cpu.decode.op21 _01454_ _01455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07520__A2 _03445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06607_ _02615_ _02928_ _02929_ _00258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_40_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07587_ _03322_ _03475_ _03483_ _00684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09326_ u_cpu.rf_ram.memory\[84\]\[2\] _04624_ _04629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06538_ u_cpu.rf_ram.memory\[47\]\[7\] _02872_ _02880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10199__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09273__A2 _04593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07284__A1 _03312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09257_ u_cpu.rf_ram.memory\[107\]\[5\] _04583_ _04589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06469_ _02669_ _02840_ _02841_ _00208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08208_ u_arbiter.i_wb_cpu_rdt\[17\] _03822_ _03833_ u_arbiter.i_wb_cpu_dbus_dat\[18\]
+ _03859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__05834__A2 _02305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09188_ _04448_ _04543_ _04550_ _01219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09025__A2 _04453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05390__S0 _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08139_ _03806_ _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08784__A1 u_arbiter.i_wb_cpu_ibus_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07587__A2 _03475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08784__B2 u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11150_ _00084_ io_in[0] u_scanchain_local.module_data_in\[62\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05598__A1 _01513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05142__S0 _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10101_ _00495_ io_in[4] u_cpu.rf_ram.memory\[52\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11081_ u_cpu.rf_ram_if.wdata1_r\[5\] io_in[4] u_cpu.rf_ram_if.wdata1_r\[4\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07339__A2 _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10032_ _00426_ io_in[4] u_cpu.rf_ram.memory\[60\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07862__C _01442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05770__A1 _01441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10934_ _01303_ io_in[4] u_cpu.rf_ram.memory\[85\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07511__A2 _03435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10865_ _01234_ io_in[4] u_cpu.rf_ram.memory\[105\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09834__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10796_ _01165_ io_in[4] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07275__A1 _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10811__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09016__A2 _04453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07027__A1 _02637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09984__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08775__A1 _03703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07578__A2 _03475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05589__A1 _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05133__S0 _01507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10961__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06250__A2 _02707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05840_ _02390_ _02399_ _00026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07750__A2 _03573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05771_ u_cpu.cpu.alu.i_rs1 _02277_ _01442_ _02346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05761__A1 _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07510_ u_cpu.rf_ram.memory\[134\]\[5\] _03435_ _03441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08490_ _03926_ _03928_ _03917_ _04093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__07502__A2 _03435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10341__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07441_ _03320_ _03395_ _03402_ _00619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07372_ _02731_ _02766_ _03364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09255__A2 _04583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09111_ u_cpu.rf_ram.memory\[101\]\[4\] _04503_ _04508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06323_ u_cpu.rf_ram.memory\[7\]\[7\] _02745_ _02753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08463__B1 _04070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10491__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09042_ _04448_ _04463_ _04470_ _01153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05816__A2 _01467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06254_ _02685_ _02707_ _02711_ _00123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09007__A2 _04436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05205_ _01602_ _01787_ _01788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05748__B u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06185_ _02628_ _02662_ _02663_ _00102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07569__A2 _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05136_ _01621_ _01719_ _01720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05124__S0 _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05067_ u_cpu.rf_ram.memory\[24\]\[1\] u_cpu.rf_ram.memory\[25\]\[1\] u_cpu.rf_ram.memory\[26\]\[1\]
+ u_cpu.rf_ram.memory\[27\]\[1\] _01508_ _01509_ _01651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09944_ _00338_ io_in[4] u_cpu.rf_ram.memory\[75\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06241__A2 _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08518__A1 _03924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08518__B2 _04000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09875_ _00269_ io_in[4] u_cpu.rf_ram.memory\[17\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09707__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09191__A1 _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08826_ u_cpu.cpu.ctrl.o_ibus_adr\[20\] _04327_ _04329_ u_cpu.cpu.ctrl.o_ibus_adr\[21\]
+ _04334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04878__I _01464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08757_ _02412_ _04293_ _04294_ _01044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_73_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05969_ u_cpu.cpu.ctrl.o_ibus_adr\[7\] _02483_ _02484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_57_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07708_ u_cpu.rf_ram.memory\[124\]\[1\] _03553_ _03555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09857__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08688_ _02392_ _03646_ _04256_ _01013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05504__A1 _01473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07639_ _03500_ _03513_ _03516_ _00703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10834__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10650_ _01023_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09309_ u_cpu.rf_ram.memory\[69\]\[4\] _04613_ _04618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08454__B1 _03988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10581_ _00954_ io_in[4] u_cpu.cpu.decode.opcode\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07009__A1 _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10984__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06480__A2 _02840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11133_ _00065_ io_in[0] u_scanchain_local.module_data_in\[45\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06232__A2 _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10214__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08509__A1 _03901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07980__A2 _03710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11064_ u_cpu.rf_ram_if.wdata0_r\[1\] io_in[4] u_cpu.rf_ram_if.wdata0_r\[0\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05991__A1 _02389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09182__A1 _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05393__B _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10015_ _00409_ io_in[4] u_cpu.rf_ram.memory\[62\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07732__A2 _03563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10364__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05743__A1 _01444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09485__A2 _04711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08532__I1 u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06299__A2 _02733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10917_ _01286_ io_in[4] u_cpu.rf_ram.memory\[59\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04929__S0 _01497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10848_ _01217_ io_in[4] u_cpu.rf_ram.memory\[99\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09237__A2 _04573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08296__I0 u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10779_ _01148_ io_in[4] u_cpu.rf_ram.memory\[96\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08996__A1 _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06471__A2 _02840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05287__C _01560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07990_ _03691_ _03720_ _03721_ _00850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07971__A2 _03710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08598__C _03972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06941_ _03106_ _03117_ _03121_ _00400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05982__A1 _02403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10707__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09173__A1 _02825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09660_ u_cpu.rf_ram.memory\[89\]\[2\] _04822_ _04825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06872_ u_cpu.rf_ram.memory\[65\]\[0\] _03079_ _03080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08611_ _02909_ u_arbiter.i_wb_cpu_rdt\[17\] _04201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05823_ _01467_ _02375_ _02385_ _00012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09591_ _04630_ _04782_ _04786_ _01386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_54_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08542_ _04138_ _04139_ _04053_ _04140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10857__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05754_ _02327_ _02328_ _02329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_54_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09476__A2 _04711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07487__A1 _03312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08473_ _03941_ _04035_ _04076_ _04077_ _04078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_51_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05685_ u_cpu.cpu.alu.i_rs1 u_cpu.cpu.alu.add_cy_r _02262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_63_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07424_ u_cpu.rf_ram.memory\[39\]\[7\] _03385_ _03393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05593__S0 _01497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07355_ _03354_ _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08987__A1 _04434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06306_ _02674_ _02742_ _02743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_137_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07286_ u_cpu.rf_ram.memory\[72\]\[3\] _03308_ _03315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09025_ u_cpu.rf_ram.memory\[95\]\[7\] _04453_ _04461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06462__A2 _02829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06237_ u_cpu.rf_ram.memory\[81\]\[4\] _02697_ _02702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10237__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06153__I _02636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06168_ _02606_ u_cpu.rf_ram_if.wdata1_r\[4\] _02649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09400__A2 _04671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05119_ _01554_ _01702_ _01607_ _01703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07411__A1 _03306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06099_ _02334_ _02588_ _02313_ _02589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07962__A2 _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09927_ _00321_ io_in[4] u_cpu.rf_ram.memory\[74\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10387__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05973__A1 u_cpu.cpu.ctrl.o_ibus_adr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09164__A1 _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09858_ _00252_ io_in[4] u_cpu.rf_ram.memory\[4\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08911__A1 _03691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07714__A2 _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08809_ _04324_ _01066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_105_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09789_ _00183_ io_in[4] u_cpu.rf_ram.memory\[46\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09467__A2 _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10702_ _01072_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08744__S _02335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06150__A1 _02606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09219__A2 _04563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05584__S0 _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11012__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10633_ _01006_ io_in[4] u_cpu.rf_ram.memory\[31\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08978__A1 _03703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10564_ _00937_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07650__A1 _02870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06453__A2 _02829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10495_ _00868_ io_in[4] u_cpu.rf_ram.memory\[11\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07953__A2 _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11116_ _00046_ io_in[0] u_arbiter.i_wb_cpu_rdt\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09155__A1 _02954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11047_ _01416_ io_in[4] u_cpu.rf_ram.memory\[89\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05716__A1 u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09458__A2 _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07469__A1 _03312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05570__C _01486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08130__A2 _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05470_ u_cpu.rf_ram.memory\[116\]\[5\] u_cpu.rf_ram.memory\[117\]\[5\] u_cpu.rf_ram.memory\[118\]\[5\]
+ u_cpu.rf_ram.memory\[119\]\[5\] _01576_ _01577_ _02050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_32_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05575__S0 _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06692__A2 _02978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07140_ u_cpu.rf_ram.memory\[53\]\[4\] _03227_ _03232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__04981__I _01504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09630__A2 _04802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07641__A1 _03502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07071_ _03110_ _03187_ _03193_ _00458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_127_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06022_ u_cpu.cpu.ctrl.o_ibus_adr\[18\] _02521_ _02526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_127_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09394__A1 _04636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08441__I0 u_arbiter.i_wb_cpu_rdt\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07944__A2 _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07973_ u_cpu.rf_ram.memory\[118\]\[1\] _03710_ _03712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05955__A1 _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09146__A1 _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09712_ _00106_ io_in[4] u_cpu.rf_ram.memory\[21\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06924_ u_cpu.rf_ram.memory\[29\]\[5\] _03100_ _03111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09643_ _04628_ _04812_ _04815_ _01409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06855_ _02881_ _03069_ _03070_ _00365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05707__A1 _01442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05806_ _02272_ u_cpu.rf_ram_if.rdata1\[4\] _02376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09574_ u_cpu.rf_ram.memory\[25\]\[4\] _04772_ _04777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06786_ _02887_ _03028_ _03031_ _00335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09449__A2 _04691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11035__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08525_ u_arbiter.i_wb_cpu_rdt\[28\] u_arbiter.i_wb_cpu_rdt\[12\] _02467_ _04125_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05737_ _02259_ _02311_ _02312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04930__A2 _01514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08121__A2 _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08456_ _03974_ _03941_ _03997_ _04050_ _03985_ _03925_ _04065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
X_05668_ _01492_ _02236_ _02245_ _02246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__05566__S0 _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07407_ _03322_ _03375_ _03383_ _00604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07880__A1 _03502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06683__A2 _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08387_ _03956_ _04007_ _04008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05599_ u_cpu.rf_ram.memory\[16\]\[7\] u_cpu.rf_ram.memory\[17\]\[7\] u_cpu.rf_ram.memory\[18\]\[7\]
+ u_cpu.rf_ram.memory\[19\]\[7\] _01508_ _01509_ _02177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_52_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07338_ u_cpu.rf_ram.memory\[70\]\[0\] _03345_ _03346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05318__S0 _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09621__A2 _04802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06435__A2 _02816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07632__A1 _02754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07269_ _02657_ _03297_ _03303_ _00546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09008_ _04450_ _04436_ _04451_ _01138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10280_ _00666_ io_in[4] u_cpu.rf_ram.memory\[132\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__04997__A2 _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06199__A1 u_cpu.cpu.immdec.imm11_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07935__A2 _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09137__A1 _02743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09688__A2 _04832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07699__A1 _03506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05174__A2 _01756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08112__A2 _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10402__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06123__A1 _02606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07871__A1 _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06674__A2 _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10616_ _00989_ io_in[4] u_cpu.cpu.immdec.imm19_12_20\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05309__S0 _01507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09612__A2 _04792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10552__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06426__A2 _02814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10547_ _00920_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08820__B1 _04329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10478_ _00851_ io_in[4] u_cpu.rf_ram.memory\[121\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09376__A1 _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07617__I _02646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05937__A1 _02403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09128__A1 _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04970_ _01494_ _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_49_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09679__A2 _04832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11058__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08351__A2 _03928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05581__B _01471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06640_ u_cpu.rf_ram.memory\[17\]\[3\] _02945_ _02949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06571_ _02637_ _02900_ _02902_ _00249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09918__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08103__A2 _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08310_ _02466_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\] _03937_ _03938_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_33_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10082__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05522_ _02094_ _02096_ _02098_ _02100_ _01541_ _02101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_09290_ _04442_ _04603_ _04607_ _01264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08241_ _03879_ _03880_ _00942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05453_ _01490_ _02023_ _02032_ _02033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__06665__A2 _02956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08172_ _03832_ _03834_ _00919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05384_ _01958_ _01960_ _01962_ _01964_ _01581_ _01965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__09603__A2 _04792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07123_ _03108_ _03217_ _03222_ _00481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06417__A2 _02805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07054_ u_cpu.rf_ram.memory\[58\]\[6\] _03177_ _03184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07090__A2 _03197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06005_ u_cpu.cpu.ctrl.o_ibus_adr\[14\] _02508_ _02512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07917__A2 _03672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09119__A1 _03037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07956_ _03699_ _03693_ _03700_ _00837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06907_ _02677_ _02803_ _03099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07887_ u_cpu.rf_ram.memory\[92\]\[7\] _03652_ _03660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06587__B _02911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08342__A2 _03961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09626_ u_cpu.rf_ram.memory\[98\]\[3\] _04802_ _04806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06838_ u_cpu.rf_ram.memory\[67\]\[1\] _03059_ _03061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10425__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06353__A1 _02681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05156__A2 _01738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09557_ _04632_ _04762_ _04767_ _01371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06769_ u_cpu.rf_ram.memory\[76\]\[3\] _03018_ _03022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08508_ _03940_ _03963_ _04109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09488_ _02259_ _02297_ _02292_ _04721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_24_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10575__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08439_ u_cpu.rf_ram.memory\[114\]\[7\] _04041_ _04049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07853__A1 _02395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06656__A2 _02956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10401_ _00774_ io_in[4] u_cpu.cpu.state.o_cnt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07605__A1 _02667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08802__B1 _04311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10332_ _00718_ io_in[4] u_cpu.rf_ram.memory\[126\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07081__A2 _03197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07865__C _02305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09358__A1 _04636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05666__B _01600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10263_ _00649_ io_in[4] u_cpu.rf_ram.memory\[134\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08030__A1 _02642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10194_ _00580_ io_in[4] u_cpu.rf_ram.memory\[70\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08581__A2 _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08333__A2 _03912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08268__I _03895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06895__A2 _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10918__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07844__A1 _03504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06647__A2 _02945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09597__A1 _04636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07072__A2 _03187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07810_ _02396_ u_cpu.cpu.state.o_cnt_r\[0\] _03613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_69_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10448__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08790_ u_cpu.cpu.ctrl.o_ibus_adr\[3\] _04309_ _04311_ u_cpu.cpu.ctrl.o_ibus_adr\[4\]
+ _04315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06583__A1 _02667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07741_ _03572_ _03573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_04953_ u_cpu.rf_ram.memory\[12\]\[0\] u_cpu.rf_ram.memory\[13\]\[0\] u_cpu.rf_ram.memory\[14\]\[0\]
+ u_cpu.rf_ram.memory\[15\]\[0\] _01530_ _01532_ _01538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_38_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09740__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08324__A2 _03912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09521__A1 _01477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07672_ u_cpu.rf_ram.memory\[126\]\[1\] _03533_ _03535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04884_ _01468_ _01470_ _01471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06335__A1 _02685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09411_ u_cpu.rf_ram.memory\[110\]\[6\] _04671_ _04678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10598__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06623_ _02889_ _02935_ _02939_ _00264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_19_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06886__A2 _03079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04897__A1 u_cpu.cpu.immdec.imm24_20\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09342_ _04638_ _04624_ _04639_ _01284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08088__A1 _03701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06554_ _02651_ _02891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09890__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05505_ u_cpu.rf_ram.memory\[28\]\[6\] u_cpu.rf_ram.memory\[29\]\[6\] u_cpu.rf_ram.memory\[30\]\[6\]
+ u_cpu.rf_ram.memory\[31\]\[6\] _01497_ _01501_ _02084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_21_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06638__A2 _02945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09273_ u_cpu.rf_ram.memory\[83\]\[4\] _04593_ _04598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06485_ _02782_ _02849_ _02850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08224_ _03868_ _03869_ _00936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05436_ _01571_ _02015_ _02016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08155_ u_arbiter.i_wb_cpu_rdt\[2\] _02924_ _03820_ _03821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05367_ u_cpu.rf_ram.memory\[100\]\[4\] u_cpu.rf_ram.memory\[101\]\[4\] u_cpu.rf_ram.memory\[102\]\[4\]
+ u_cpu.rf_ram.memory\[103\]\[4\] _01551_ _01524_ _01948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_101_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07106_ u_cpu.rf_ram.memory\[55\]\[5\] _03207_ _03213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08086_ _03699_ _03770_ _03774_ _00893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07063__A2 _03187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05298_ u_cpu.rf_ram.memory\[92\]\[3\] u_cpu.rf_ram.memory\[93\]\[3\] u_cpu.rf_ram.memory\[94\]\[3\]
+ u_cpu.rf_ram.memory\[95\]\[3\] _01562_ _01563_ _01880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_134_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05486__B _01519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07037_ _02662_ _03167_ _03174_ _00443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06810__A2 _03039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08012__A1 _02642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06023__B1 _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08563__A2 _04009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08988_ _02636_ _04438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07939_ u_cpu.rf_ram.memory\[117\]\[6\] _03682_ _03689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09512__A1 u_cpu.cpu.genblk3.csr.mstatus_mie vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10950_ _01319_ io_in[4] u_cpu.rf_ram.memory\[86\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05129__A2 _01712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06326__A1 _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09609_ _02685_ _04792_ _04796_ _01394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_10881_ _01250_ io_in[4] u_cpu.rf_ram.memory\[107\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06877__A2 _03079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07826__A1 _03504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06629__A2 _02935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08752__S _02335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09579__A1 _04636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08251__A1 _03691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07054__A2 _03177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10315_ _00701_ io_in[4] u_cpu.rf_ram.memory\[128\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06801__A2 _03039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10246_ _00632_ io_in[4] u_cpu.rf_ram.memory\[136\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09763__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08554__A2 _03998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10177_ _00563_ io_in[4] u_cpu.rf_ram.memory\[73\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06565__A1 _02897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10740__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06868__A2 _03069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04879__A1 u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10890__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06270_ _02681_ _02719_ _02721_ _00129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07293__A2 _03308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10120__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05221_ u_cpu.rf_ram.memory\[68\]\[2\] u_cpu.rf_ram.memory\[69\]\[2\] u_cpu.rf_ram.memory\[70\]\[2\]
+ u_cpu.rf_ram.memory\[71\]\[2\] _01507_ _01605_ _01804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_128_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08242__A1 u_arbiter.i_wb_cpu_rdt\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05152_ _01473_ _01686_ _01735_ _00001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07045__A2 _03177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05083_ u_cpu.rf_ram.memory\[36\]\[1\] u_cpu.rf_ram.memory\[37\]\[1\] u_cpu.rf_ram.memory\[38\]\[1\]
+ u_cpu.rf_ram.memory\[39\]\[1\] _01544_ _01545_ _01667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09960_ _00354_ io_in[4] u_cpu.rf_ram.memory\[68\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10270__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08911_ _03691_ _04381_ _04382_ _01110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09891_ _00285_ io_in[4] u_cpu.rf_ram.memory\[119\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08842_ u_cpu.cpu.ctrl.o_ibus_adr\[28\] _04327_ _04329_ u_cpu.cpu.ctrl.o_ibus_adr\[29\]
+ _04342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06556__A1 _02891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08773_ _03701_ _04299_ _04304_ _01050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05985_ _02403_ u_scanchain_local.module_data_in\[47\] _02478_ u_arbiter.i_wb_cpu_dbus_adr\[10\]
+ _02497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_85_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07724_ u_cpu.rf_ram.memory\[123\]\[0\] _03563_ _03564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04936_ _01503_ _01511_ _01515_ _01520_ _01486_ _01521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_84_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06859__A2 _03069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07655_ _03498_ _03523_ _03525_ _00710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04867_ u_cpu.cpu.decode.op26 _01454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06606_ u_cpu.rf_ram_if.rcnt\[0\] u_cpu.rf_ram_if.rcnt\[2\] u_cpu.rf_ram_if.rcnt\[1\]
+ _02929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_07586_ u_cpu.rf_ram.memory\[130\]\[7\] _03475_ _03483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09325_ _02641_ _04628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06537_ _02691_ _02872_ _02879_ _00238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07808__A1 u_cpu.cpu.state.o_cnt_r\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09256_ _04444_ _04583_ _04588_ _01249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06468_ u_cpu.rf_ram.memory\[41\]\[0\] _02840_ _02841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08481__A1 _04069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07284__A2 _03308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05295__A1 _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08207_ u_arbiter.i_wb_cpu_dbus_dat\[17\] _03835_ _03858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05419_ u_cpu.rf_ram.memory\[24\]\[5\] u_cpu.rf_ram.memory\[25\]\[5\] u_cpu.rf_ram.memory\[26\]\[5\]
+ u_cpu.rf_ram.memory\[27\]\[5\] _01508_ _01509_ _01999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09187_ u_cpu.rf_ram.memory\[99\]\[6\] _04543_ _04550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06399_ _02687_ _02794_ _02799_ _00180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10613__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05390__S1 _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08138_ u_arbiter.i_wb_cpu_ack _02397_ _03806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__07036__A2 _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05047__A1 _01492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09786__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08784__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08069_ u_cpu.rf_ram.memory\[122\]\[4\] _03760_ _03765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05142__S1 _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10100_ _00494_ io_in[4] u_cpu.rf_ram.memory\[52\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11080_ u_cpu.rf_ram_if.wdata1_r\[4\] io_in[4] u_cpu.rf_ram_if.wdata1_r\[3\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10763__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10031_ _00425_ io_in[4] u_cpu.rf_ram.memory\[60\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06547__A1 _02885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11119__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10933_ _01302_ io_in[4] u_cpu.rf_ram.memory\[85\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10864_ _01233_ io_in[4] u_cpu.rf_ram.memory\[105\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10143__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10795_ _01164_ io_in[4] u_cpu.rf_ram.memory\[28\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07275__A2 _02954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05286__A1 _01566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05676__I3 u_cpu.rf_ram.memory\[139\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10293__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07027__A2 _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08775__A2 _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05589__A2 _02167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06786__A1 _02887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05133__S1 _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10229_ _00615_ io_in[4] u_cpu.rf_ram.memory\[137\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05770_ _01441_ _02344_ _02345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05761__A2 _02335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07440_ u_cpu.rf_ram.memory\[137\]\[6\] _03395_ _03402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06710__A1 _02881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07371_ _03322_ _03355_ _03363_ _00588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09110_ _04442_ _04503_ _04507_ _01184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10636__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06322_ _02662_ _02745_ _02752_ _00150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_31_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07266__A2 _03297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08463__A1 u_cpu.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05277__A1 _01490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09041_ u_cpu.rf_ram.memory\[96\]\[6\] _04463_ _04470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06253_ u_cpu.rf_ram.memory\[18\]\[3\] _02707_ _02711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05204_ u_cpu.rf_ram.memory\[112\]\[2\] u_cpu.rf_ram.memory\[113\]\[2\] u_cpu.rf_ram.memory\[114\]\[2\]
+ u_cpu.rf_ram.memory\[115\]\[2\] _01572_ _01545_ _01787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_129_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07018__A2 _03157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06184_ u_cpu.rf_ram.memory\[82\]\[6\] _02628_ _02663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05029__A1 _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10786__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08766__A2 _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05135_ u_cpu.rf_ram.memory\[72\]\[1\] u_cpu.rf_ram.memory\[73\]\[1\] u_cpu.rf_ram.memory\[74\]\[1\]
+ u_cpu.rf_ram.memory\[75\]\[1\] _01522_ _01622_ _01719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_144_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05124__S1 _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05066_ _01493_ _01649_ _01650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09943_ _00337_ io_in[4] u_cpu.rf_ram.memory\[75\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08518__A2 _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10016__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06529__A1 _02683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09874_ _00268_ io_in[4] u_cpu.rf_ram.memory\[16\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09191__A2 _02870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08825_ _04333_ _01073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05201__A1 _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05968_ u_cpu.cpu.ctrl.o_ibus_adr\[6\] u_cpu.cpu.ctrl.o_ibus_adr\[5\] _02476_ _02483_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08756_ _02355_ _04293_ _04294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10166__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07707_ _03494_ _03553_ _03554_ _00733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_04919_ u_cpu.cpu.csr_imm u_cpu.rf_ram_if.rtrig0 _01453_ _01461_ _01504_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_54_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05899_ u_arbiter.i_wb_cpu_rdt\[20\] u_arbiter.i_wb_cpu_dbus_dat\[17\] _02431_ _02436_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08687_ u_cpu.cpu.alu.cmp_r _02392_ _04256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04894__I _01480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07638_ u_cpu.rf_ram.memory\[128\]\[2\] _03513_ _03516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05060__S0 _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07569_ _03322_ _03465_ _03473_ _00676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_16_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09308_ _04442_ _04613_ _04617_ _01272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10580_ _00953_ io_in[4] u_cpu.rf_ram.memory\[113\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08454__A1 _03899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08454__B2 _03925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09239_ u_cpu.rf_ram.memory\[106\]\[5\] _04573_ _04579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07009__A2 _03157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05658__C _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08757__A2 _04293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06768__A1 _02887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11132_ _00064_ io_in[0] u_scanchain_local.module_data_in\[44\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05440__A1 _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11063_ _01431_ io_in[4] u_cpu.cpu.state.ibus_cyc vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10014_ _00408_ io_in[4] u_cpu.rf_ram.memory\[62\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09182__A2 _04543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10509__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07193__A1 _02647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05743__A2 _02265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09801__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11091__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10659__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10916_ _01285_ io_in[4] u_cpu.rf_ram.memory\[59\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07496__A2 _03425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04929__S1 _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05051__S0 _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10847_ _01216_ io_in[4] u_cpu.rf_ram.memory\[99\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09951__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08445__A1 _03935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07248__A2 _03287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10778_ _01147_ io_in[4] u_cpu.rf_ram.memory\[96\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08996__A2 _04436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07799__A3 _03605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10039__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07420__A2 _03385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05431__A1 _01528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06940_ u_cpu.rf_ram.memory\[63\]\[3\] _03117_ _03121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09173__A2 _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10189__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06871_ _03078_ _03079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_41_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07184__A1 _02731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08920__A2 _04381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08610_ u_cpu.cpu.immdec.imm19_12_20\[6\] _04165_ _04200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05822_ u_cpu.rf_ram_if.rdata0\[5\] _01467_ _02385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09590_ u_cpu.rf_ram.memory\[24\]\[3\] _04782_ _04786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06931__A1 _03114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05290__S0 _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08541_ _03932_ _03918_ _04128_ _04139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05753_ u_cpu.cpu.decode.opcode\[1\] _02328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_36_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08472_ _04034_ _04077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08684__A1 _03705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07487__A2 _03425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05684_ u_arbiter.i_wb_cpu_dbus_we u_cpu.cpu.bufreg.i_sh_signed _02260_ _01445_ _02261_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_78_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07423_ _03320_ _03385_ _03392_ _00611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05042__S0 _01522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05593__S1 _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07354_ _02870_ _02976_ _03354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08436__A1 _03703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06305_ _02616_ _02671_ _02742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08987__A2 _04436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07285_ _02646_ _03314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09024_ _04448_ _04453_ _04460_ _01145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06236_ _02685_ _02697_ _02701_ _00115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06167_ _02628_ _02647_ _02648_ _00099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05118_ u_cpu.rf_ram.memory\[116\]\[1\] u_cpu.rf_ram.memory\[117\]\[1\] u_cpu.rf_ram.memory\[118\]\[1\]
+ u_cpu.rf_ram.memory\[119\]\[1\] _01576_ _01577_ _01702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_85_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07411__A2 _03385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06098_ _02587_ _02329_ _02305_ _02588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_78_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05422__A1 _01513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05049_ _01522_ _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09926_ _00320_ io_in[4] u_cpu.rf_ram.memory\[74\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09164__A2 _04533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09824__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09857_ _00251_ io_in[4] u_cpu.rf_ram.memory\[4\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07175__A1 _02647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08911__A2 _04381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08808_ u_cpu.cpu.ctrl.o_ibus_adr\[12\] _04309_ _04311_ u_cpu.cpu.ctrl.o_ibus_adr\[13\]
+ _04324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08297__S _02464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06922__A1 _03108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09788_ _00182_ io_in[4] u_cpu.rf_ram.memory\[46\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10801__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05281__S0 _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08739_ _04282_ _01038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09974__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07478__A2 _03415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05033__S0 _01507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10701_ _01071_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10951__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05584__S1 _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10632_ _01005_ io_in[4] u_cpu.rf_ram.memory\[31\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08978__A2 _04425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05669__B _01471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10563_ _00936_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06989__A1 _03098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07650__A2 _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08760__S _04293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10494_ _00867_ io_in[4] u_cpu.rf_ram.memory\[11\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07402__A2 _03375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10331__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05949__C1 _02398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05413__A1 _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11115_ _00045_ io_in[0] u_arbiter.i_wb_cpu_rdt\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09155__A2 _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11046_ _01415_ io_in[4] u_cpu.rf_ram.memory\[89\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07166__A1 _02731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08902__A2 _04371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10481__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06913__A1 _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05272__S0 _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07469__A2 _03415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08666__A1 _03705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05575__S1 _01563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08418__A1 _03969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08969__A2 _04425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09091__A1 u_arbiter.i_wb_cpu_rdt\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07070_ u_cpu.rf_ram.memory\[57\]\[5\] _03187_ _03193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07641__A2 _03513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06021_ _02525_ _00076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_126_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09394__A2 _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09847__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08441__I1 u_arbiter.i_wb_cpu_rdt\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05404__A1 _01492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07972_ _03691_ _03710_ _03711_ _00842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10824__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09146__A2 _04523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09711_ _00105_ io_in[4] u_cpu.rf_ram.memory\[21\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06923_ _02656_ _03110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07157__A1 _03106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09997__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09642_ u_cpu.rf_ram.memory\[100\]\[2\] _04812_ _04815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06854_ u_cpu.rf_ram.memory\[66\]\[0\] _03069_ _03070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05707__A2 _01439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05263__S0 _01551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05805_ _02273_ u_cpu.rf_ram.rdata\[4\] _02375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09573_ _04630_ _04772_ _04776_ _01378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06785_ u_cpu.rf_ram.memory\[75\]\[2\] _03028_ _03031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10974__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06380__A2 _02784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08524_ _03896_ _04101_ _04124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05736_ _01445_ _02265_ _02310_ _01444_ _02311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_36_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05667_ _02238_ _02240_ _02242_ _02244_ _01541_ _02245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_08455_ _04053_ _04062_ _04063_ _03901_ _04064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_24_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05566__S1 _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10204__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07406_ u_cpu.rf_ram.memory\[138\]\[7\] _03375_ _03383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08386_ _03974_ _03904_ _03969_ _04006_ _04007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__08409__A1 _03910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07880__A2 _03652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05598_ _01513_ _02175_ _02176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07337_ _03344_ _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05318__S1 _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07268_ u_cpu.rf_ram.memory\[13\]\[5\] _03297_ _03303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07632__A2 _02976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10354__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05643__A1 _01566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09007_ u_cpu.rf_ram.memory\[94\]\[7\] _04436_ _04451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06219_ _02689_ _02679_ _02690_ _00109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07199_ _02662_ _03257_ _03264_ _00515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09385__A2 _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06199__A2 u_cpu.cpu.immdec.imm11_7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08593__B1 _04183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09137__A2 _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09909_ _00303_ io_in[4] u_cpu.rf_ram.memory\[139\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07148__A1 _02717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07699__A2 _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05254__S0 _01523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08648__A1 _02263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05006__S0 _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06123__A2 _02303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07871__A2 _02814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10615_ _00988_ io_in[4] u_cpu.cpu.immdec.imm19_12_20\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05309__S1 _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10546_ _00919_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05634__A1 _01548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10477_ _00850_ io_in[4] u_cpu.rf_ram.memory\[121\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10847__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09376__A2 _04651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07387__A1 _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09128__A2 _04513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07139__A1 _03106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10997__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11029_ _01398_ io_in[4] u_cpu.rf_ram.memory\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08887__A1 _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05245__S0 _01497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06362__A2 _02770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10227__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06570_ u_cpu.rf_ram.memory\[4\]\[1\] _02900_ _02902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08639__A1 _02305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05521_ _01513_ _02099_ _01482_ _02100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_75_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07311__A1 _03316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08240_ u_arbiter.i_wb_cpu_rdt\[28\] _03807_ _03829_ u_arbiter.i_wb_cpu_dbus_dat\[29\]
+ _03880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__04992__I _01498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05452_ _02025_ _02027_ _02029_ _02031_ _01581_ _02032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_20_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07862__A2 _02334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10377__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08171_ u_arbiter.i_wb_cpu_dbus_dat\[5\] _03808_ _03833_ _02922_ _03834_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05383_ _01554_ _01963_ _01607_ _01964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07122_ u_cpu.rf_ram.memory\[54\]\[4\] _03217_ _03222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05102__B _01685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05625__A1 _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07053_ _03110_ _03177_ _03183_ _00450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_12_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06004_ _02463_ _02510_ _02511_ _00073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09367__A2 _04651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05928__A2 _02403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09119__A2 _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06050__A1 _02461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11002__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07955_ u_cpu.rf_ram.memory\[120\]\[3\] _03693_ _03700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08327__B1 _03915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06906_ _02631_ _03098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07886_ _03508_ _03652_ _03659_ _00808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05236__S0 _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09625_ _04628_ _04802_ _04805_ _01401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06837_ _02881_ _03059_ _03060_ _00357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05491__C _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06353__A2 _02770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09556_ u_cpu.rf_ram.memory\[26\]\[4\] _04762_ _04767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11152__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06159__I _02641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06768_ _02887_ _03018_ _03021_ _00327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08507_ _03944_ _03975_ _04093_ _04108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_93_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05719_ u_cpu.cpu.genblk3.csr.mcause3_0\[0\] _02295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_102_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09487_ _02263_ _02303_ _04720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06699_ u_cpu.rf_ram.memory\[129\]\[4\] _02978_ _02983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08438_ _03705_ _04041_ _04048_ _00971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05164__I0 u_cpu.rf_ram.memory\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05864__A1 _02416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09055__A1 _04438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08369_ _03935_ _03984_ _03985_ _03986_ _03991_ _03992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_109_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10400_ _00773_ io_in[4] u_cpu.cpu.state.stage_two_req vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07605__A2 _03485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05616__A1 _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10331_ _00717_ io_in[4] u_cpu.rf_ram.memory\[126\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10262_ _00648_ io_in[4] u_cpu.rf_ram.memory\[134\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09358__A2 _04641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07369__A1 _03320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08030__A2 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10193_ _00579_ io_in[4] u_cpu.rf_ram.memory\[70\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05919__A2 _02403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06041__A1 _02456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06592__A2 u_arbiter.i_wb_cpu_dbus_dat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08869__A1 _03705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09530__A2 _04752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07541__A1 _03312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09294__A1 _04446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08097__A2 _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07844__A2 _03626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09046__A1 _04141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09597__A2 _04782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05607__A1 _01528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10529_ _00902_ io_in[4] u_cpu.rf_ram.memory\[116\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06280__A1 _02691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09349__A2 _04641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11025__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08021__A2 _03730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06032__A1 _02389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05466__S0 _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06583__A2 _02900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04987__I _01495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04952_ _01528_ _01536_ _01537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07740_ _02782_ _03037_ _03572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09521__A2 _02301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07671_ _03494_ _03533_ _03534_ _00717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_04883_ u_cpu.cpu.immdec.imm24_20\[4\] _01469_ _01470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06335__A2 _02756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09410_ _04634_ _04671_ _04677_ _01314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06622_ u_cpu.rf_ram.memory\[16\]\[3\] _02935_ _02939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09341_ u_cpu.rf_ram.memory\[84\]\[7\] _04624_ _04639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06553_ _02889_ _02883_ _02890_ _00243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08088__A2 _03770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06099__A1 _02334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05504_ _01473_ _02034_ _02083_ _00005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06484_ _02742_ _02779_ _02849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09272_ _04442_ _04593_ _04597_ _01256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07835__A2 _03626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05846__A1 _02400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08223_ u_arbiter.i_wb_cpu_rdt\[22\] _03807_ _03829_ u_arbiter.i_wb_cpu_dbus_dat\[23\]
+ _03869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05435_ u_cpu.rf_ram.memory\[36\]\[5\] u_cpu.rf_ram.memory\[37\]\[5\] u_cpu.rf_ram.memory\[38\]\[5\]
+ u_cpu.rf_ram.memory\[39\]\[5\] _01544_ _01545_ _02015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_14_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09588__A2 _04782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08154_ _03816_ _03818_ _02924_ _03819_ _03820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05366_ _01492_ _01918_ _01927_ _01946_ _01947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_14_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07599__A1 _02652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08796__B1 _04311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07105_ _03108_ _03207_ _03212_ _00473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08085_ u_cpu.rf_ram.memory\[115\]\[3\] _03770_ _03774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08260__A2 _03885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05297_ _01490_ _01869_ _01878_ _01879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_07036_ u_cpu.rf_ram.memory\[5\]\[6\] _03167_ _03174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08012__A2 _03730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05457__S0 _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06023__A1 _02402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08987_ _04434_ _04436_ _04437_ _01131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06574__A2 _02900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07771__A1 _03506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07938_ _03506_ _03682_ _03688_ _00831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10542__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07869_ u_cpu.cpu.state.init_done _03611_ _03650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07523__A1 _03312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06326__A2 _02754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09608_ u_cpu.rf_ram.memory\[0\]\[3\] _04792_ _04796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05007__B _01558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10880_ _01249_ io_in[4] u_cpu.rf_ram.memory\[107\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09539_ _04632_ _04752_ _04757_ _01363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08079__A2 _03770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09276__A1 _04446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10692__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07826__A2 _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05837__A1 _02396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09579__A2 _04772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11048__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05677__B _01534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08251__A2 _03885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06262__A1 _02693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10314_ _00700_ io_in[4] u_cpu.rf_ram.memory\[22\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09908__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09200__A1 _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08003__A2 _03720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10245_ _00631_ io_in[4] u_cpu.rf_ram.memory\[136\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10072__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05448__S0 _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10176_ _00562_ io_in[4] u_cpu.rf_ram.memory\[73\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06565__A2 _02883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06317__A2 _02745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04879__A2 _01452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05620__S0 _01496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07817__A2 _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08490__A2 _03928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06096__A4 _02585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05220_ _01621_ _01802_ _01803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05151_ _01725_ _01734_ _01735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08242__A2 _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10415__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05082_ _01659_ _01661_ _01663_ _01665_ _01541_ _01666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_100_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08910_ u_cpu.rf_ram.memory\[93\]\[0\] _04381_ _04382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09890_ _00284_ io_in[4] u_cpu.rf_ram.memory\[40\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06005__A1 u_cpu.cpu.ctrl.o_ibus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05439__S0 _01551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08841_ _04341_ _01081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10565__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06556__A2 _02883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07753__A1 _03506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08772_ u_cpu.rf_ram.memory\[30\]\[4\] _04299_ _04304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05984_ u_cpu.cpu.ctrl.o_ibus_adr\[10\] _02493_ _02496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_84_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07723_ _03562_ _03563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_04935_ _01506_ _01516_ _01519_ _01520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07505__A1 _03312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07654_ u_cpu.rf_ram.memory\[127\]\[1\] _03523_ _03525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_04866_ _01440_ _01452_ _01453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_92_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06605_ u_cpu.rf_ram_if.rcnt\[0\] _02928_ _00257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05611__S0 _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09258__A1 _04446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07585_ _03320_ _03475_ _03482_ _00683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09324_ _04626_ _04624_ _04627_ _01278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05382__I3 u_cpu.rf_ram.memory\[119\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06536_ u_cpu.rf_ram.memory\[47\]\[6\] _02872_ _02879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07808__A2 _03611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05819__A1 _01467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09255_ u_cpu.rf_ram.memory\[107\]\[4\] _04583_ _04588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06467_ _02839_ _02840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08481__A2 _04083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05295__A2 _01876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06492__A1 _02683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08206_ _03856_ _03857_ _00930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05418_ _01493_ _01997_ _01998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09186_ _04446_ _04543_ _04549_ _01218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06398_ u_cpu.rf_ram.memory\[46\]\[4\] _02794_ _02799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08137_ u_arbiter.i_wb_cpu_dbus_dat\[1\] _02915_ _02924_ _03805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05497__B _01534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05349_ u_cpu.rf_ram.memory\[32\]\[4\] u_cpu.rf_ram.memory\[33\]\[4\] u_cpu.rf_ram.memory\[34\]\[4\]
+ u_cpu.rf_ram.memory\[35\]\[4\] _01495_ _01499_ _01930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09430__A1 _04636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08233__A2 _03874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10095__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06244__A1 _02693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08068_ _03699_ _03760_ _03764_ _00885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10908__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07992__A1 _03695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06795__A2 _03028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07019_ _03112_ _03157_ _03164_ _00435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10030_ _00424_ io_in[4] u_cpu.rf_ram.memory\[60\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06547__A2 _02883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10932_ _01301_ io_in[4] u_cpu.rf_ram.memory\[85\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05602__S0 _01523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10863_ _01232_ io_in[4] u_cpu.rf_ram.memory\[105\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06347__I _02767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10794_ _01163_ io_in[4] u_cpu.rf_ram.memory\[28\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10438__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06483__A1 _02693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09730__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10588__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06786__A2 _03028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08511__B _03938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09880__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10228_ _00614_ io_in[4] u_cpu.rf_ram.memory\[137\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07735__A1 _03506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06538__A2 _02872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10159_ _00545_ io_in[4] u_cpu.rf_ram.memory\[13\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09488__A1 _02259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08160__B2 _03802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06710__A2 _02988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07370_ u_cpu.rf_ram.memory\[143\]\[7\] _03355_ _03363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06321_ u_cpu.rf_ram.memory\[7\]\[6\] _02745_ _02752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08463__A2 _04069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09040_ _04446_ _04463_ _04469_ _01152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06252_ _02683_ _02707_ _02710_ _00122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05277__A2 _01849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05203_ _01597_ _01785_ _01600_ _01786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06183_ _02661_ _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09412__A1 _04636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05110__B _01558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05134_ _01617_ _01717_ _01519_ _01718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06777__A2 _03018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07974__A1 _03695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05065_ u_cpu.rf_ram.memory\[28\]\[1\] u_cpu.rf_ram.memory\[29\]\[1\] u_cpu.rf_ram.memory\[30\]\[1\]
+ u_cpu.rf_ram.memory\[31\]\[1\] _01497_ _01501_ _01649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09942_ _00336_ io_in[4] u_cpu.rf_ram.memory\[75\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09517__B _02396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05985__B1 _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09873_ _00267_ io_in[4] u_cpu.rf_ram.memory\[16\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06529__A2 _02872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08824_ u_cpu.cpu.ctrl.o_ibus_adr\[19\] _04327_ _04329_ u_cpu.cpu.ctrl.o_ibus_adr\[20\]
+ _04333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08755_ _02596_ _02914_ _04292_ _04293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05967_ _02456_ _02481_ _02482_ _00064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_73_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07706_ u_cpu.rf_ram.memory\[124\]\[0\] _03553_ _03554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04918_ _01493_ _01502_ _01503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08686_ _03707_ _04247_ _04255_ _01012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05898_ _02435_ _00040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08151__A1 u_arbiter.i_wb_cpu_dbus_dat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07637_ _03498_ _03513_ _03515_ _00702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04849_ _01436_ u_cpu.rf_ram_if.rcnt\[2\] u_cpu.rf_ram_if.rcnt\[1\] _01437_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_53_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06701__A2 _02978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05060__S1 _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07568_ u_cpu.rf_ram.memory\[131\]\[7\] _03465_ _03473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09307_ u_cpu.rf_ram.memory\[69\]\[3\] _04613_ _04617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06519_ u_cpu.rf_ram.memory\[48\]\[7\] _02861_ _02869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09753__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09651__A1 _04636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08454__A2 _03975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07499_ _03434_ _03435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_16_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09238_ _04444_ _04573_ _04578_ _01241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10730__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09169_ u_cpu.rf_ram.memory\[104\]\[6\] _04533_ _04540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06116__B _02392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07965__A1 _03705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06768__A2 _03018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11131_ _00063_ io_in[0] u_scanchain_local.module_data_in\[43\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10880__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05440__A2 _02019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11062_ _01430_ io_in[4] u_cpu.rf_ram.memory\[23\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07717__A1 _03506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10013_ _00407_ io_in[4] u_cpu.rf_ram.memory\[62\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07193__A2 _03257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10110__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06940__A2 _03117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10915_ _01284_ io_in[4] u_cpu.rf_ram.memory\[84\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10260__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05051__S1 _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10846_ _01215_ io_in[4] u_cpu.rf_ram.memory\[99\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10777_ _01146_ io_in[4] u_cpu.rf_ram.memory\[95\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08445__A2 _03974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06456__A1 _02685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07956__A1 _03699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06759__A2 _03008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05431__A2 _02010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06540__I _02631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06870_ _02695_ _02768_ _03078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08381__A1 _03965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07184__A2 _02870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05821_ _01467_ _02373_ _02384_ _00011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06931__A2 _03100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08540_ _03922_ _03923_ _04004_ _04137_ _03998_ _04138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_78_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05290__S1 _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05752_ _02265_ _02327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__04942__A1 _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08467__I u_cpu.cpu.immdec.imm24_20\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10603__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08133__A1 _02259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08471_ _03970_ _03971_ _04022_ _04076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09776__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05683_ _01441_ u_cpu.cpu.bne_or_bge _02260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_36_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08684__A2 _04247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07422_ u_cpu.rf_ram.memory\[39\]\[6\] _03385_ _03392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05042__S1 _01622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10753__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07353_ _03322_ _03345_ _03353_ _00580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09633__A1 _04636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08436__A2 _04041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08416__B _03915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06447__A1 _02825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06304_ _02667_ _02733_ _02741_ _00143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07284_ _03312_ _03308_ _03313_ _00551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06998__A2 _03147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09023_ u_cpu.rf_ram.memory\[95\]\[6\] _04453_ _04460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06235_ u_cpu.rf_ram.memory\[81\]\[3\] _02697_ _02701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11109__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06166_ u_cpu.rf_ram.memory\[82\]\[3\] _02628_ _02648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07947__A1 _03691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05117_ _01602_ _01700_ _01701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06097_ _02265_ u_cpu.cpu.decode.opcode\[1\] _02587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08151__B _02915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05048_ _01610_ _01632_ _01471_ _01633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05422__A2 _02001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09925_ _00319_ io_in[4] u_cpu.rf_ram.memory\[74\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10133__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09856_ _00250_ io_in[4] u_cpu.rf_ram.memory\[4\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07175__A2 _03247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08372__A1 _03965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08807_ _04323_ _01065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_100_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09787_ _00181_ io_in[4] u_cpu.rf_ram.memory\[46\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06999_ _03110_ _03147_ _03153_ _00426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06922__A2 _03100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10283__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05281__S1 _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08738_ u_arbiter.i_wb_cpu_dbus_adr\[26\] u_arbiter.i_wb_cpu_dbus_adr\[27\] _02335_
+ _04282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08124__A1 _03701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08669_ _02677_ _02870_ _04246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08675__A2 _04247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10700_ _01070_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05033__S1 _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10631_ _01004_ io_in[4] u_cpu.rf_ram.memory\[32\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08427__A2 _04041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10562_ _00935_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06989__A2 _03147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05110__A1 _01566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10493_ _00866_ io_in[4] u_cpu.rf_ram.memory\[11\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07938__A1 _03506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05949__B1 _02463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05949__C2 u_arbiter.i_wb_cpu_dbus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11114_ _00044_ io_in[0] u_arbiter.i_wb_cpu_rdt\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05413__A2 _01993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06610__A1 _02912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11045_ _01414_ io_in[4] u_cpu.rf_ram.memory\[100\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10626__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08363__A1 _03914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07166__A2 _02838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05905__S _02431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09799__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06913__A2 _03100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05716__A3 _02291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05272__S1 _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10776__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08666__A2 _04237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06677__A1 _02887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10829_ _01198_ io_in[4] u_cpu.rf_ram.memory\[103\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09615__A1 _02691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10006__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06429__A1 _02669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05579__C _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09091__A2 _04485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05101__A1 _01490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06020_ _02389_ u_scanchain_local.module_data_in\[54\] _02524_ _02525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10156__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05404__A2 _01975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06601__A1 _02313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07971_ u_cpu.rf_ram.memory\[118\]\[0\] _03710_ _03711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09710_ _00104_ io_in[4] u_cpu.rf_ram.memory\[21\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06922_ _03108_ _03100_ _03109_ _00393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08354__A1 _02466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07157__A2 _03237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09641_ _04626_ _04812_ _04814_ _01408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06853_ _03068_ _03069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06904__A2 _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05804_ _02272_ _02373_ _02374_ _00017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_82_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09572_ u_cpu.rf_ram.memory\[25\]\[3\] _04772_ _04776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05263__S1 _01524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06784_ _02885_ _03028_ _03030_ _00334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08106__A1 _03701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08523_ _03966_ _04121_ _04122_ _04123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_64_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05735_ _02285_ _02309_ _02260_ _02310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08657__A2 _04237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06668__A1 _02897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08454_ _03899_ _03975_ _03988_ _03925_ _03938_ _04063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_05666_ _01617_ _02243_ _01600_ _02244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_24_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07405_ _03320_ _03375_ _03382_ _00603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08385_ _04000_ _03918_ _03930_ _03945_ _04005_ _04006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__09606__A1 u_cpu.rf_ram.memory\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05597_ u_cpu.rf_ram.memory\[20\]\[7\] u_cpu.rf_ram.memory\[21\]\[7\] u_cpu.rf_ram.memory\[22\]\[7\]
+ u_cpu.rf_ram.memory\[23\]\[7\] _01530_ _01532_ _02175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_104_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07336_ _02768_ _03037_ _03344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07093__A1 _03114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07267_ _02652_ _03297_ _03302_ _00545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_87_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09006_ _02666_ _04450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_139_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06218_ u_cpu.rf_ram.memory\[21\]\[5\] _02679_ _02690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07198_ u_cpu.rf_ram.memory\[15\]\[6\] _03257_ _03264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11081__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06149_ _02628_ _02632_ _02633_ _00096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10649__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08593__A1 _01439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07396__A2 _03375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09941__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09908_ _00302_ io_in[4] u_cpu.rf_ram.memory\[139\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08345__A1 _03909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07148__A2 _02827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09839_ _00233_ io_in[4] u_cpu.rf_ram.memory\[47\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10799__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08896__A2 _04371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05254__S1 _01525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08648__A2 _02598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10029__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05006__S1 _01531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07320__A2 _03335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10614_ _00987_ io_in[4] u_cpu.cpu.immdec.imm19_12_20\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10179__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10545_ _00918_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08820__A2 _04327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06831__A1 _02895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10476_ _00849_ io_in[4] u_cpu.rf_ram.memory\[118\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08584__A1 _03910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07387__A2 _03365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05398__A1 _01617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08336__A1 _03906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07139__A2 _03227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11028_ _01397_ io_in[4] u_cpu.rf_ram.memory\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08887__A2 _04361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05245__S1 _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05520_ u_cpu.rf_ram.memory\[12\]\[6\] u_cpu.rf_ram.memory\[13\]\[6\] u_cpu.rf_ram.memory\[14\]\[6\]
+ u_cpu.rf_ram.memory\[15\]\[6\] _01530_ _01532_ _02099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_17_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07311__A2 _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05451_ _01597_ _02030_ _01579_ _02031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_75_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08170_ _03829_ _03833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05382_ u_cpu.rf_ram.memory\[116\]\[4\] u_cpu.rf_ram.memory\[117\]\[4\] u_cpu.rf_ram.memory\[118\]\[4\]
+ u_cpu.rf_ram.memory\[119\]\[4\] _01576_ _01577_ _01963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09814__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09064__A2 _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07121_ _03106_ _03217_ _03221_ _00480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07075__A1 _03114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05625__A2 _02202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07052_ u_cpu.rf_ram.memory\[58\]\[5\] _03177_ _03183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06003_ _02402_ u_scanchain_local.module_data_in\[51\] _02478_ u_arbiter.i_wb_cpu_dbus_adr\[14\]
+ _02511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_133_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09964__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07378__A2 _03365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05389__A1 _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10941__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07954_ _02646_ _03699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08327__A1 _03944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08327__B2 _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06905_ _02897_ _03089_ _03097_ _00388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07885_ u_cpu.rf_ram.memory\[92\]\[6\] _03652_ _03659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08878__A2 _04361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09624_ u_cpu.rf_ram.memory\[98\]\[2\] _04802_ _04805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06836_ u_cpu.rf_ram.memory\[67\]\[0\] _03059_ _03060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05236__S1 _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07550__A2 _03455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09555_ _04630_ _04762_ _04766_ _01370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06767_ u_cpu.rf_ram.memory\[76\]\[2\] _03018_ _03021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05561__A1 _01490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08506_ _04067_ _04107_ _00980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05718_ u_cpu.cpu.state.o_cnt_r\[3\] _02290_ _02292_ _02293_ _02294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_09486_ _04638_ _04711_ _04719_ _01348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06698_ _02889_ _02978_ _02982_ _00296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07302__A2 _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10321__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08437_ u_cpu.rf_ram.memory\[114\]\[6\] _04041_ _04048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05649_ _01490_ _02217_ _02226_ _02227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__05864__A2 _02389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08368_ _03915_ _03990_ _03991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09055__A2 _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07319_ _03334_ _03335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08299_ _02464_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[8\] _03927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08802__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10471__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10330_ _00716_ io_in[4] u_cpu.rf_ram.memory\[127\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06813__A1 _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05616__A2 _02193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10261_ _00647_ io_in[4] u_cpu.rf_ram.memory\[134\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08566__A1 _04160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07369__A2 _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08566__B2 _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10192_ _00578_ io_in[4] u_cpu.rf_ram.memory\[70\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06592__A3 u_arbiter.i_wb_cpu_dbus_dat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08869__A2 _04351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07541__A2 _03455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11087__CLKN io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09837__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09294__A2 _04603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10814__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05203__B _01600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07057__A1 _03114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09987__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10528_ _00901_ io_in[4] u_cpu.rf_ram.memory\[116\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10964__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06280__A2 _02719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10459_ _00832_ io_in[4] u_cpu.rf_ram.memory\[117\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08557__A1 _03925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05466__S1 _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08309__A1 _02466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07780__A2 _03593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04951_ u_cpu.rf_ram.memory\[8\]\[0\] u_cpu.rf_ram.memory\[9\]\[0\] u_cpu.rf_ram.memory\[10\]\[0\]
+ u_cpu.rf_ram.memory\[11\]\[0\] _01523_ _01525_ _01536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_38_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05791__A1 _02363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11166__I io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07670_ u_cpu.rf_ram.memory\[126\]\[0\] _03533_ _03534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04882_ _01438_ _01452_ _01469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_65_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07532__A2 _03445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10344__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06621_ _02887_ _02935_ _02938_ _00263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09340_ _02666_ _04638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06552_ u_cpu.rf_ram.memory\[50\]\[3\] _02883_ _02890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09285__A2 _04603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04936__C _01486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05503_ _02073_ _02082_ _02083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07296__A1 _03320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09271_ u_cpu.rf_ram.memory\[83\]\[3\] _04593_ _04597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06483_ _02693_ _02840_ _02848_ _00215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10494__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08222_ u_arbiter.i_wb_cpu_dbus_dat\[22\] _03808_ _03868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05846__A2 _02398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05434_ _02007_ _02009_ _02011_ _02013_ _01541_ _02014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_14_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09037__A2 _04463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08153_ u_arbiter.i_wb_cpu_dbus_dat\[2\] _03812_ _03819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08245__B1 _03833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05365_ _01490_ _01936_ _01945_ _01946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_88_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07599__A2 _03485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07104_ u_cpu.rf_ram.memory\[55\]\[4\] _03207_ _03212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08796__B2 u_cpu.cpu.ctrl.o_ibus_adr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08084_ _03697_ _03770_ _03773_ _00892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05296_ _01871_ _01873_ _01875_ _01877_ _01581_ _01878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_49_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07035_ _02657_ _03167_ _03173_ _00442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06271__A2 _02719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07220__A1 _02803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05457__S1 _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08986_ u_cpu.rf_ram.memory\[94\]\[0\] _04436_ _04437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07771__A2 _03583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07937_ u_cpu.rf_ram.memory\[117\]\[5\] _03682_ _03688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05909__I0 u_arbiter.i_wb_cpu_rdt\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07868_ _03649_ _00800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07523__A2 _03445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06819_ _02881_ _03049_ _03050_ _00349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_3_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09607_ _02683_ _04792_ _04795_ _01393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_113_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07799_ _02395_ _03604_ _03605_ _00774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_43_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09538_ u_cpu.rf_ram.memory\[27\]\[4\] _04752_ _04757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10837__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09276__A2 _04593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07287__A1 _03314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09469_ _02626_ _02954_ _04710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06119__B _02604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05023__B _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07039__A1 _02667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10987__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04862__B u_cpu.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10313_ _00699_ io_in[4] u_cpu.rf_ram.memory\[22\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06262__A2 _02707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10217__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08539__A1 _03923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10244_ _00630_ io_in[4] u_cpu.rf_ram.memory\[136\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09200__A2 _04553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07211__A1 _03106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05448__S1 _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10175_ _00561_ io_in[4] u_cpu.rf_ram.memory\[73\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07762__A2 _03583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10367__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05773__A1 u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08496__S _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07514__A2 _03435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05913__S _02431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05620__S1 _01594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09267__A2 _04593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07278__A1 _03306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09019__A2 _04453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08490__A3 _03917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05150_ _01727_ _01729_ _01731_ _01733_ _01466_ _01734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__06253__A2 _02707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05081_ _01513_ _01664_ _01482_ _01665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11142__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08840_ u_cpu.cpu.ctrl.o_ibus_adr\[27\] _04327_ _04329_ u_cpu.cpu.ctrl.o_ibus_adr\[28\]
+ _04341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07202__A1 _02766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05439__S1 _01524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08950__A1 u_cpu.cpu.immdec.imm11_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07753__A2 _03573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08771_ _03699_ _04299_ _04303_ _01049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05983_ _02493_ _02494_ _02495_ _00067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07722_ _02849_ _02965_ _03562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04934_ _01518_ _01519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07505__A2 _03435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07653_ _03494_ _03523_ _03524_ _00709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04865_ _01447_ _01449_ _01451_ _01452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06604_ _02912_ _02927_ _02928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07584_ u_cpu.rf_ram.memory\[130\]\[6\] _03475_ _03482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05611__S1 _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09258__A2 _04583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09323_ u_cpu.rf_ram.memory\[84\]\[1\] _04624_ _04627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07269__A1 _02657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06535_ _02689_ _02872_ _02878_ _00237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09254_ _04442_ _04583_ _04587_ _01248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05819__A2 _02371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06466_ _02782_ _02838_ _02839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08205_ u_arbiter.i_wb_cpu_rdt\[16\] _03822_ _03833_ u_arbiter.i_wb_cpu_dbus_dat\[17\]
+ _03857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05417_ u_cpu.rf_ram.memory\[28\]\[5\] u_cpu.rf_ram.memory\[29\]\[5\] u_cpu.rf_ram.memory\[30\]\[5\]
+ u_cpu.rf_ram.memory\[31\]\[5\] _01497_ _01501_ _01997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09185_ u_cpu.rf_ram.memory\[99\]\[5\] _04543_ _04549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06492__A2 _02851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06397_ _02685_ _02794_ _02798_ _00179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08154__B _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08769__A1 _03697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08136_ _03802_ _03803_ _03804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05348_ _01543_ _01928_ _01929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09430__A2 _04681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05047__A3 _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07441__A1 _03320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06244__A2 _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08067_ u_cpu.rf_ram.memory\[122\]\[3\] _03760_ _03764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05279_ u_cpu.rf_ram.memory\[100\]\[3\] u_cpu.rf_ram.memory\[101\]\[3\] u_cpu.rf_ram.memory\[102\]\[3\]
+ u_cpu.rf_ram.memory\[103\]\[3\] _01551_ _01573_ _01861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_88_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07992__A2 _03720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07018_ u_cpu.rf_ram.memory\[19\]\[6\] _03157_ _03164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09194__A1 _04434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08601__C _03969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08941__A1 _03986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07744__A2 _03573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08969_ u_cpu.rf_ram.memory\[97\]\[1\] _04425_ _04427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10931_ _01300_ io_in[4] u_cpu.rf_ram.memory\[10\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10862_ _01231_ io_in[4] u_cpu.rf_ram.memory\[105\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05602__S1 _01525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09249__A2 _04583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06180__A1 _02606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11015__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10793_ _01162_ io_in[4] u_cpu.rf_ram.memory\[28\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06483__A2 _02840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05118__S0 _01576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09421__A2 _04681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06235__A2 _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07983__A2 _03710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10227_ _00613_ io_in[4] u_cpu.rf_ram.memory\[137\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07735__A2 _03563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08932__A1 _03928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10158_ _00544_ io_in[4] u_cpu.rf_ram.memory\[13\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05746__A1 _02263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10089_ _00483_ io_in[4] u_cpu.rf_ram.memory\[54\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08999__A1 _04444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06320_ _02657_ _02745_ _02751_ _00149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09660__A2 _04822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06251_ u_cpu.rf_ram.memory\[18\]\[2\] _02707_ _02710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06474__A2 _02840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05277__A3 _01858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07671__A1 _03494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05202_ u_cpu.rf_ram.memory\[120\]\[2\] u_cpu.rf_ram.memory\[121\]\[2\] u_cpu.rf_ram.memory\[122\]\[2\]
+ u_cpu.rf_ram.memory\[123\]\[2\] _01598_ _01556_ _01785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_102_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05109__S0 _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06182_ _02660_ _02661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09412__A2 _04671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10532__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07423__A1 _03320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05133_ u_cpu.rf_ram.memory\[68\]\[1\] u_cpu.rf_ram.memory\[69\]\[1\] u_cpu.rf_ram.memory\[70\]\[1\]
+ u_cpu.rf_ram.memory\[71\]\[1\] _01507_ _01605_ _01717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_85_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07974__A2 _03710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05064_ _01473_ _01584_ _01648_ _00000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09941_ _00335_ io_in[4] u_cpu.rf_ram.memory\[75\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05985__A1 _02403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09176__A1 _04434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08421__C _03955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09872_ _00266_ io_in[4] u_cpu.rf_ram.memory\[16\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10682__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07726__A2 _03563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08923__A1 _03705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08823_ _04332_ _01072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05737__A1 _02259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08754_ u_cpu.cpu.state.o_cnt_r\[1\] u_cpu.cpu.state.o_cnt_r\[0\] _02292_ _02914_
+ _04292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05966_ _02418_ u_scanchain_local.module_data_in\[43\] _02398_ u_arbiter.i_wb_cpu_dbus_adr\[6\]
+ _02482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_38_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09479__A2 _04711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07705_ _03552_ _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11038__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04917_ u_cpu.rf_ram.memory\[28\]\[0\] u_cpu.rf_ram.memory\[29\]\[0\] u_cpu.rf_ram.memory\[30\]\[0\]
+ u_cpu.rf_ram.memory\[31\]\[0\] _01497_ _01501_ _01502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_26_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08685_ u_cpu.rf_ram.memory\[31\]\[7\] _04247_ _04255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05897_ u_arbiter.i_wb_cpu_rdt\[19\] u_arbiter.i_wb_cpu_dbus_dat\[16\] _02431_ _02435_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08151__A2 u_arbiter.i_wb_cpu_dbus_dat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07636_ u_cpu.rf_ram.memory\[128\]\[1\] _03513_ _03515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04848_ u_cpu.rf_ram_if.rcnt\[0\] _01436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06162__A1 _02606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07567_ _03320_ _03465_ _03472_ _00675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10062__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09306_ _04440_ _04613_ _04616_ _01271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06518_ _02691_ _02861_ _02868_ _00230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_70_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07498_ _02976_ _03037_ _03434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09651__A2 _04812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09237_ u_cpu.rf_ram.memory\[106\]\[4\] _04573_ _04578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06449_ u_cpu.rf_ram.memory\[51\]\[0\] _02829_ _02830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07279__I _02636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05301__B _01600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06183__I _02661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09168_ _04446_ _04533_ _04539_ _01210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09403__A2 _04671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08119_ u_cpu.rf_ram.memory\[33\]\[2\] _03790_ _03793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09099_ u_arbiter.i_wb_cpu_rdt\[31\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\]
+ _02910_ _04501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_107_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07965__A2 _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11130_ _00062_ io_in[0] u_scanchain_local.module_data_in\[42\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06911__I _02636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05976__A1 _02456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05520__S0 _01530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11061_ _01429_ io_in[4] u_cpu.rf_ram.memory\[23\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07717__A2 _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10012_ _00406_ io_in[4] u_cpu.rf_ram.memory\[62\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05728__A1 u_arbiter.i_wb_cpu_ibus_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10405__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10914_ _01283_ io_in[4] u_cpu.rf_ram.memory\[84\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10845_ _01214_ io_in[4] u_cpu.rf_ram.memory\[99\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10776_ _01145_ io_in[4] u_cpu.rf_ram.memory\[95\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09642__A2 _04812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10555__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07653__A1 _03494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06456__A2 _02829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07405__A1 _03320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07956__A2 _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05967__A1 _02456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05511__S0 _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09158__A1 _04434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07708__A2 _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08905__A1 _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08381__A2 _03972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05820_ u_cpu.rf_ram_if.rdata0\[4\] _01467_ _02384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05751_ _01445_ u_arbiter.i_wb_cpu_dbus_we _02325_ _01457_ _02326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__04942__A2 _01526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10085__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09330__A1 _04630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08470_ u_arbiter.i_wb_cpu_rdt\[23\] u_arbiter.i_wb_cpu_rdt\[7\] _02466_ _04075_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05682_ _02258_ _02259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_62_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07421_ _03318_ _03385_ _03391_ _00610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_78_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07892__A1 _03494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06695__A2 _02978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07352_ u_cpu.rf_ram.memory\[70\]\[7\] _03345_ _03353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09633__A2 _04802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06303_ u_cpu.rf_ram.memory\[1\]\[7\] _02733_ _02741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06447__A2 _02827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07283_ u_cpu.rf_ram.memory\[72\]\[2\] _03308_ _03313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09022_ _04446_ _04453_ _04459_ _01144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06234_ _02683_ _02697_ _02700_ _00114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09397__A1 _02766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06165_ _02646_ _02647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07947__A2 _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05116_ u_cpu.rf_ram.memory\[112\]\[1\] u_cpu.rf_ram.memory\[113\]\[1\] u_cpu.rf_ram.memory\[114\]\[1\]
+ u_cpu.rf_ram.memory\[115\]\[1\] _01544_ _01545_ _01700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__05958__A1 _02456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05775__C _02336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06096_ u_cpu.cpu.alu.i_rs1 u_cpu.cpu.bufreg.c_r _02584_ _02585_ _02586_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_49_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05047_ _01492_ _01620_ _01631_ _01632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_09924_ _00318_ io_in[4] u_cpu.rf_ram.memory\[74\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09855_ _00249_ io_in[4] u_cpu.rf_ram.memory\[4\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08372__A2 _03961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08806_ u_cpu.cpu.ctrl.o_ibus_adr\[11\] _04309_ _04311_ u_cpu.cpu.ctrl.o_ibus_adr\[12\]
+ _04323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__05791__B _01460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10428__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09786_ _00180_ io_in[4] u_cpu.rf_ram.memory\[46\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06998_ u_cpu.rf_ram.memory\[60\]\[5\] _03147_ _03153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06383__A1 _02689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05949_ _02389_ u_scanchain_local.module_data_in\[39\] _02463_ _02468_ _02398_ u_arbiter.i_wb_cpu_dbus_adr\[2\]
+ _02469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
X_08737_ _04281_ _01037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09720__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09321__A1 _04622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08124__A2 _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08594__S _02466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06135__A1 u_cpu.cpu.immdec.imm11_7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08668_ _03707_ _04237_ _04245_ _01004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10578__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07619_ _03502_ _03496_ _03503_ _00696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06686__A2 _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08599_ _03932_ _03998_ _04190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10630_ _01003_ io_in[4] u_cpu.rf_ram.memory\[32\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06906__I _02631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09870__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09624__A2 _04802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06438__A2 _02816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10561_ _00934_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07635__A1 _03494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08832__B1 _04329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10492_ _00865_ io_in[4] u_cpu.rf_ram.memory\[8\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09388__A1 _04630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07938__A2 _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05949__A1 _02389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11113_ _00043_ io_in[0] u_arbiter.i_wb_cpu_rdt\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06610__A2 _02927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11044_ _01413_ io_in[4] u_cpu.rf_ram.memory\[100\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08363__A2 _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08115__A2 _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09312__A1 _04446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07874__A1 _03494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06677__A2 _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10828_ _01197_ io_in[4] u_cpu.rf_ram.memory\[103\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09615__A2 _04792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06429__A2 _02816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10759_ _01128_ io_in[4] u_cpu.rf_ram.memory\[97\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05101__A2 _01675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09379__A1 _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07929__A2 _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04860__A1 _01443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06551__I _02646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06062__B1 _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07970_ _03709_ _03710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05404__A3 _01984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06921_ u_cpu.rf_ram.memory\[29\]\[4\] _03100_ _03109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09743__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09551__A1 _04626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09640_ u_cpu.rf_ram.memory\[100\]\[1\] _04812_ _04814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06852_ _02619_ _02768_ _03068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06365__A1 _02693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05803_ _02272_ u_cpu.rf_ram_if.rdata1\[3\] _02374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09571_ _04628_ _04772_ _04775_ _01377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06783_ u_cpu.rf_ram.memory\[75\]\[1\] _03028_ _03030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10720__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08106__A2 _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08522_ _03924_ _03910_ _04051_ _04122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_05734_ _01442_ _02309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_70_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06117__A1 u_cpu.cpu.immdec.imm11_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09893__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08453_ _04057_ _04059_ _04061_ _04062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_35_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05665_ u_cpu.rf_ram.memory\[76\]\[7\] u_cpu.rf_ram.memory\[77\]\[7\] u_cpu.rf_ram.memory\[78\]\[7\]
+ u_cpu.rf_ram.memory\[79\]\[7\] _01529_ _01500_ _02243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07865__A1 _02265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06668__A2 _02956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07404_ u_cpu.rf_ram.memory\[138\]\[6\] _03375_ _03382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10870__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08384_ _03970_ _04004_ _04005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05596_ _01506_ _02173_ _01481_ _02174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_91_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09606__A2 _04792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07335_ _03322_ _03335_ _03343_ _00572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08290__A1 _03906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07266_ u_cpu.rf_ram.memory\[13\]\[4\] _03297_ _03302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07093__A2 _03197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10100__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09005_ _04448_ _04436_ _04449_ _01137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06217_ _02656_ _02689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06840__A2 _03059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07197_ _02657_ _03257_ _03263_ _00514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06148_ u_cpu.rf_ram.memory\[82\]\[0\] _02628_ _02633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08593__A2 _04165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06199__A4 _02622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06079_ _02402_ u_scanchain_local.module_data_in\[65\] _02478_ u_arbiter.i_wb_cpu_dbus_adr\[28\]
+ _02573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10250__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09907_ _00301_ io_in[4] u_cpu.rf_ram.memory\[139\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08345__A2 _03917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09838_ _00232_ io_in[4] u_cpu.rf_ram.memory\[47\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09769_ _00163_ io_in[4] u_cpu.rf_ram.memory\[78\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06659__A2 _02956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07856__A1 u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__04865__B _01451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08337__B _03962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10613_ _00986_ io_in[4] u_cpu.cpu.immdec.imm19_12_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10544_ _00917_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07084__A2 _03197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08281__A1 _03906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05095__A1 _01566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10475_ _00848_ io_in[4] u_cpu.rf_ram.memory\[118\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06831__A2 _03049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09081__I0 u_arbiter.i_wb_cpu_rdt\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09766__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08584__A2 _03985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06595__A1 _02915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10743__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08336__A2 _03947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09533__A1 _04626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11027_ _01396_ io_in[4] u_cpu.rf_ram.memory\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06898__A2 _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10893__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05570__A2 _02144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05858__B1 _02413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05450_ u_cpu.rf_ram.memory\[48\]\[5\] u_cpu.rf_ram.memory\[49\]\[5\] u_cpu.rf_ram.memory\[50\]\[5\]
+ u_cpu.rf_ram.memory\[51\]\[5\] _01576_ _01577_ _02030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_61_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10123__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05381_ _01602_ _01961_ _01962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07120_ u_cpu.rf_ram.memory\[54\]\[3\] _03217_ _03221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07075__A2 _03187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05086__A1 _01548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07051_ _03108_ _03177_ _03182_ _00449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06822__A2 _03049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10273__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06002_ u_cpu.cpu.ctrl.o_ibus_adr\[14\] _02508_ _02510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_133_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06035__B1 _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06586__A1 _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07953_ _03697_ _03693_ _03698_ _00836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08327__A2 _03912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09524__A1 u_cpu.cpu.ctrl.i_iscomp vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06904_ u_cpu.rf_ram.memory\[64\]\[7\] _03089_ _03097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07884_ _03506_ _03652_ _03658_ _00807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09623_ _04626_ _04802_ _04804_ _01400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06835_ _03058_ _03059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09554_ u_cpu.rf_ram.memory\[26\]\[3\] _04762_ _04766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06766_ _02885_ _03018_ _03020_ _00326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_93_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05561__A2 _02130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08505_ u_cpu.cpu.immdec.imm30_25\[1\] _04104_ _04106_ u_cpu.cpu.immdec.imm30_25\[2\]
+ _04107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05717_ u_cpu.cpu.decode.op26 _01447_ _02293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07838__A1 _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09485_ u_cpu.rf_ram.memory\[88\]\[7\] _04711_ _04719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06697_ u_cpu.rf_ram.memory\[129\]\[3\] _02978_ _02982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08436_ _03703_ _04041_ _04047_ _00970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05648_ _02219_ _02221_ _02223_ _02225_ _01581_ _02226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_12_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06510__A1 _02683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08367_ _03970_ _03987_ _03989_ _03990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05579_ _02151_ _02153_ _02155_ _02157_ _01541_ _02158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__10616__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07318_ _02743_ _02768_ _03334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08263__A1 _03705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07066__A2 _03187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08298_ _03922_ _03923_ _03924_ _03925_ _03926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XANTENNA__05077__A1 _01528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09789__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07249_ _03108_ _03287_ _03292_ _00537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06813__A2 _03039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05872__I0 u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10260_ _00646_ io_in[4] u_cpu.rf_ram.memory\[134\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10766__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10191_ _00577_ io_in[4] u_cpu.rf_ram.memory\[70\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06577__A1 _02652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08318__A2 _03944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09515__A1 u_cpu.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06592__A4 u_arbiter.i_wb_cpu_dbus_dat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06329__A1 _02669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05001__A1 _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10146__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10296__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07057__A2 _03177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05068__A1 _01506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08514__C _03966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10527_ _00900_ io_in[4] u_cpu.rf_ram.memory\[116\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06804__A2 _03039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10458_ _00831_ io_in[4] u_cpu.rf_ram.memory\[117\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08557__A2 _03948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10389_ _00762_ io_in[4] u_cpu.rf_ram.memory\[37\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08309__A2 _02411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05240__A1 _01473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04950_ _01528_ _01533_ _01534_ _01535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_78_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04881_ u_cpu.cpu.immdec.imm19_12_20\[8\] _01467_ _01468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08190__B1 _03833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06620_ u_cpu.rf_ram.memory\[16\]\[2\] _02935_ _02938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06740__A1 _02895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11071__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06551_ _02646_ _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05502_ _02075_ _02077_ _02079_ _02081_ _01466_ _02082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_09270_ _04440_ _04593_ _04596_ _01255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10639__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08493__A1 _03901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08692__S _04257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07296__A2 _03308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06482_ u_cpu.rf_ram.memory\[41\]\[7\] _02840_ _02848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08221_ _03866_ _03867_ _00935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05433_ _01513_ _02012_ _01482_ _02013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09931__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08152_ _03802_ _03817_ _03818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07048__A2 _03177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05364_ _01938_ _01940_ _01942_ _01944_ _01581_ _01945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05059__A1 _01465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10789__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07103_ _03106_ _03207_ _03211_ _00472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08083_ u_cpu.rf_ram.memory\[115\]\[2\] _03770_ _03773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08796__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05295_ _01554_ _01876_ _01607_ _01877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07034_ u_cpu.rf_ram.memory\[5\]\[5\] _03167_ _03173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10019__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06559__A1 _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07220__A2 _02976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08985_ _04435_ _04436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_76_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05231__A1 _01465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07936_ _03504_ _03682_ _03687_ _00830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05782__A2 _02356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10169__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07867_ u_cpu.cpu.mem_bytecnt\[1\] u_cpu.cpu.state.o_cnt\[2\] _02291_ _00780_ _03649_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_56_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08181__B1 _03833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09606_ u_cpu.rf_ram.memory\[0\]\[2\] _04792_ _04795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06818_ u_cpu.rf_ram.memory\[68\]\[0\] _03049_ _03050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07798_ u_cpu.cpu.state.o_cnt_r\[3\] u_cpu.cpu.state.o_cnt\[2\] _03605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_43_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09537_ _04630_ _04752_ _04756_ _01362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06749_ u_cpu.rf_ram.memory\[74\]\[2\] _03008_ _03011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06186__I u_cpu.rf_ram_if.wdata1_r\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09468_ _04638_ _04701_ _04709_ _01340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_12_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07287__A2 _03308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06119__C _02598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08419_ _04035_ _04036_ _04037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09399_ u_cpu.rf_ram.memory\[110\]\[0\] _04671_ _04672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07039__A2 _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06914__I _02641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06798__A1 _02731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10312_ _00698_ io_in[4] u_cpu.rf_ram.memory\[22\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08539__A2 _03935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10243_ _00629_ io_in[4] u_cpu.rf_ram.memory\[136\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07211__A2 _03267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10174_ _00560_ io_in[4] u_cpu.rf_ram.memory\[73\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05222__A1 _01617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09804__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11094__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06722__A1 _02895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09954__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08475__A1 _03906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07278__A2 _03308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05289__A1 _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10931__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08778__A2 _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05080_ u_cpu.rf_ram.memory\[12\]\[1\] u_cpu.rf_ram.memory\[13\]\[1\] u_cpu.rf_ram.memory\[14\]\[1\]
+ u_cpu.rf_ram.memory\[15\]\[1\] _01530_ _01532_ _01664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07450__A2 _03405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07202__A2 _02976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10311__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05213__A1 _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08770_ u_cpu.rf_ram.memory\[30\]\[3\] _04299_ _04303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05982_ _02403_ u_scanchain_local.module_data_in\[46\] _02478_ u_arbiter.i_wb_cpu_dbus_adr\[9\]
+ _02495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_97_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05764__A2 _02330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06961__A1 _03108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07721_ _03510_ _03553_ _03561_ _00740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_04933_ _01517_ _01518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10461__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07652_ u_cpu.rf_ram.memory\[127\]\[0\] _03523_ _03524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04864_ _01450_ _01446_ u_cpu.cpu.genblk3.csr.o_new_irq u_cpu.cpu.state.genblk1.misalign_trap_sync_r
+ _01451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_53_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06713__A1 u_cpu.rf_ram.memory\[139\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06603_ _02305_ _02925_ _02926_ _02927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07583_ _03318_ _03475_ _03481_ _00682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06534_ u_cpu.rf_ram.memory\[47\]\[5\] _02872_ _02878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09322_ _02636_ _04626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08466__A1 _04029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07269__A2 _03297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09253_ u_cpu.rf_ram.memory\[107\]\[3\] _04583_ _04587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06465_ _02672_ _02779_ _02838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08204_ u_arbiter.i_wb_cpu_dbus_dat\[16\] _03835_ _03856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05416_ _01473_ _01947_ _01996_ _00004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09184_ _04444_ _04543_ _04548_ _01217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06396_ u_cpu.rf_ram.memory\[46\]\[3\] _02794_ _02798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08769__A2 _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08135_ u_arbiter.i_wb_cpu_dbus_dat\[0\] _02915_ _03803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05347_ u_cpu.rf_ram.memory\[36\]\[4\] u_cpu.rf_ram.memory\[37\]\[4\] u_cpu.rf_ram.memory\[38\]\[4\]
+ u_cpu.rf_ram.memory\[39\]\[4\] _01544_ _01545_ _01928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_107_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08066_ _03697_ _03760_ _03763_ _00884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07441__A2 _03395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05278_ _01492_ _01831_ _01840_ _01859_ _01860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_134_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07017_ _03110_ _03157_ _03163_ _00434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09827__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09194__A2 _04553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08968_ _03691_ _04425_ _04426_ _01123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10804__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07919_ u_cpu.rf_ram.memory\[34\]\[5\] _03672_ _03678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08899_ _02647_ _04371_ _04375_ _01105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_84_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09977__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10930_ _01299_ io_in[4] u_cpu.rf_ram.memory\[10\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06704__A1 _02895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10861_ _01230_ io_in[4] u_cpu.rf_ram.memory\[105\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10954__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05034__B _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08457__A1 _03910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10792_ _01161_ io_in[4] u_cpu.rf_ram.memory\[28\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07680__A2 _03533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05691__A1 u_arbiter.i_wb_cpu_dbus_we vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05118__S1 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07432__A2 _03395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10334__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05994__A2 _02499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09185__A2 _04543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10226_ _00612_ io_in[4] u_cpu.rf_ram.memory\[39\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10157_ _00543_ io_in[4] u_cpu.rf_ram.memory\[13\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10484__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06943__A1 _03108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05597__I2 u_cpu.rf_ram.memory\[22\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05924__S _02431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10088_ _00482_ io_in[4] u_cpu.rf_ram.memory\[54\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09488__A3 _02292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05054__S0 _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08448__A1 _04052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08999__A2 _04436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06250_ _02681_ _02707_ _02709_ _00121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06554__I _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07671__A2 _03533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05201_ _01543_ _01783_ _01784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06181_ _02611_ u_cpu.rf_ram_if.wdata0_r\[6\] _02659_ _02660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_117_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05109__S1 _01531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05132_ _01621_ _01715_ _01716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08620__A1 _04164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07423__A2 _03385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05434__A1 _02007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05063_ _01633_ _01647_ _01648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09940_ _00334_ io_in[4] u_cpu.rf_ram.memory\[75\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10827__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09176__A2 _04543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09871_ _00265_ io_in[4] u_cpu.rf_ram.memory\[16\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07187__A1 _02632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08923__A2 _04381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08822_ u_cpu.cpu.ctrl.o_ibus_adr\[18\] _04327_ _04329_ u_cpu.cpu.ctrl.o_ibus_adr\[19\]
+ _04332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05119__B _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08753_ _04291_ _01043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05965_ u_cpu.cpu.ctrl.o_ibus_adr\[6\] _02480_ _02481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10977__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07704_ _02814_ _02965_ _03552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04916_ _01500_ _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08684_ _03705_ _04247_ _04254_ _01011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05896_ _02434_ _00039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08151__A3 u_arbiter.i_wb_cpu_dbus_dat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07635_ _03494_ _03513_ _03514_ _00701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10207__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07566_ u_cpu.rf_ram.memory\[131\]\[6\] _03465_ _03472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09305_ u_cpu.rf_ram.memory\[69\]\[2\] _04613_ _04616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06517_ u_cpu.rf_ram.memory\[48\]\[6\] _02861_ _02868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07497_ _03322_ _03425_ _03433_ _00644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_16_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07111__A1 _03114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09236_ _04442_ _04573_ _04577_ _01240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07662__A2 _03523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06448_ _02828_ _02829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10357__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05673__A1 _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09167_ u_cpu.rf_ram.memory\[104\]\[5\] _04533_ _04539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06379_ _02685_ _02784_ _02788_ _00171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08118_ _03695_ _03790_ _03792_ _00907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08611__A1 _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07414__A2 _03385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09098_ _04500_ _01179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_79_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08049_ u_cpu.rf_ram.memory\[112\]\[3\] _03750_ _03754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05520__S1 _01532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09167__A2 _04533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11060_ _01428_ io_in[4] u_cpu.rf_ram.memory\[23\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10011_ _00405_ io_in[4] u_cpu.rf_ram.memory\[62\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08914__A2 _04381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05029__B _01600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06925__A1 _03110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05728__A2 _02303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08678__A1 _03699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10913_ _01282_ io_in[4] u_cpu.rf_ram.memory\[84\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11132__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10844_ _01213_ io_in[4] u_cpu.rf_ram.memory\[99\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10775_ _01144_ io_in[4] u_cpu.rf_ram.memory\[95\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07653__A2 _03523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08850__A1 _01451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05664__A1 _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08602__A1 _03928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07405__A2 _03375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05416__A1 _01473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05511__S1 _01509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09158__A2 _04533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07169__A1 _02632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08366__B1 _03988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10209_ _00595_ io_in[4] u_cpu.rf_ram.memory\[14\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08905__A2 _04371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06916__A1 _03104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06392__A2 _02794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05750_ u_cpu.cpu.decode.co_ebreak _02325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08669__A1 _02677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09330__A2 _04624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05681_ u_cpu.cpu.state.o_cnt_r\[1\] u_cpu.cpu.state.o_cnt_r\[0\] u_cpu.cpu.state.o_cnt_r\[3\]
+ u_cpu.cpu.state.o_cnt_r\[2\] _02258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_36_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06144__A2 _02606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07341__A1 _03310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07420_ u_cpu.rf_ram.memory\[39\]\[5\] _03385_ _03391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07892__A2 _03662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07351_ _03320_ _03345_ _03352_ _00579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06302_ _02662_ _02733_ _02740_ _00142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05402__B _01481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07282_ _02641_ _03312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07644__A2 _03513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09021_ u_cpu.rf_ram.memory\[95\]\[5\] _04453_ _04459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05655__A1 _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06233_ u_cpu.rf_ram.memory\[81\]\[2\] _02697_ _02700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09397__A2 _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06164_ _02645_ _02646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05407__A1 _01465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05115_ _01597_ _01698_ _01600_ _01699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_105_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06095_ _01445_ _02327_ _02585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09149__A2 _04523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05046_ _01624_ _01626_ _01628_ _01630_ _01541_ _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_09923_ _00317_ io_in[4] u_cpu.rf_ram.memory\[74\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11005__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09854_ _00248_ io_in[4] u_cpu.rf_ram.memory\[4\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06907__A1 _02677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08805_ _04322_ _01064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_100_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09785_ _00179_ io_in[4] u_cpu.rf_ram.memory\[46\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06997_ _03108_ _03147_ _03152_ _00425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06383__A2 _02784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11155__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08736_ u_arbiter.i_wb_cpu_dbus_adr\[25\] u_arbiter.i_wb_cpu_dbus_adr\[26\] _02335_
+ _04281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_73_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05948_ _02467_ u_cpu.cpu.ctrl.o_ibus_adr\[2\] _02468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05018__S0 _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09321__A2 _04624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08667_ u_cpu.rf_ram.memory\[32\]\[7\] _04237_ _04245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05879_ _02425_ _00030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06135__A2 _02608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07618_ u_cpu.rf_ram.memory\[22\]\[3\] _03496_ _03503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07883__A2 _03652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08598_ _03940_ _03929_ _03975_ _03972_ _04189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_26_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07549_ _03320_ _03455_ _03462_ _00667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10560_ _00933_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07635__A2 _03513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09219_ u_cpu.rf_ram.memory\[105\]\[4\] _04563_ _04568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10491_ _00864_ io_in[4] u_cpu.rf_ram.memory\[8\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08623__B _03910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09388__A2 _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07399__A1 _03314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11112_ _00042_ io_in[0] u_arbiter.i_wb_cpu_rdt\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11043_ _01412_ io_in[4] u_cpu.rf_ram.memory\[100\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08899__A1 _02647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09560__A2 _04762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06374__A2 _02784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09312__A2 _04613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10522__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07323__A1 _03310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07874__A2 _03652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10827_ _01196_ io_in[4] u_cpu.rf_ram.memory\[102\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05222__B _01519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10672__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10758_ _01127_ io_in[4] u_cpu.rf_ram.memory\[97\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10689_ _01059_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05101__A3 _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09379__A2 _02675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11028__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08051__A2 _03750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06062__A1 _02402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05496__S0 _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06920_ _02651_ _03108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10052__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09551__A2 _04762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06851_ _02897_ _03059_ _03067_ _00364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06365__A2 _02770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05802_ _02273_ u_cpu.rf_ram.rdata\[3\] _02373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09570_ u_cpu.rf_ram.memory\[25\]\[2\] _04772_ _04775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06782_ _02881_ _03028_ _03029_ _00333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08521_ _04118_ _04120_ _04053_ _04121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09303__A2 _04613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05733_ _01445_ _02303_ _02307_ _02308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_24_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06117__A2 u_cpu.cpu.immdec.imm11_7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08452_ _04060_ _04061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05664_ _01602_ _02241_ _02242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07403_ _03318_ _03375_ _03381_ _00602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05595_ u_cpu.rf_ram.memory\[24\]\[7\] u_cpu.rf_ram.memory\[25\]\[7\] u_cpu.rf_ram.memory\[26\]\[7\]
+ u_cpu.rf_ram.memory\[27\]\[7\] _01522_ _01622_ _02173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08383_ _03942_ _03971_ _04004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09067__A1 _04450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07334_ u_cpu.rf_ram.memory\[71\]\[7\] _03335_ _03343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07265_ _02647_ _03297_ _03301_ _00544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08290__A2 _03917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09004_ u_cpu.rf_ram.memory\[94\]\[6\] _04436_ _04449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06216_ _02687_ _02679_ _02688_ _00108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07196_ u_cpu.rf_ram.memory\[15\]\[5\] _03257_ _03263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_3_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06147_ _02631_ _02632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06053__A1 _02389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05487__S0 _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06078_ _02456_ _02571_ _02572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05800__A1 _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05029_ _01597_ _01613_ _01600_ _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_59_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09906_ _00300_ io_in[4] u_cpu.rf_ram.memory\[129\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09542__A2 _04752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09837_ _00231_ io_in[4] u_cpu.rf_ram.memory\[48\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10545__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06356__A2 _02770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06189__I _02666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09768_ _00162_ io_in[4] u_cpu.rf_ram.memory\[78\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08719_ _04272_ _01028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09699_ u_cpu.rf_ram_if.rcnt\[0\] u_cpu.rf_ram_if.rcnt\[1\] _04846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07305__A1 _03310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10695__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06917__I _02646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10612_ _00985_ io_in[4] u_cpu.cpu.immdec.imm7 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10543_ _00916_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08281__A2 _03908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06292__A1 _02637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10474_ _00847_ io_in[4] u_cpu.rf_ram.memory\[118\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10075__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09230__A1 _04434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08033__A2 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05478__S0 _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06601__B _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09533__A2 _04752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11026_ _01395_ io_in[4] u_cpu.rf_ram.memory\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05217__B _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05650__S0 _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07847__A2 _03626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05858__A1 _02411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09049__A1 _02395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05380_ u_cpu.rf_ram.memory\[112\]\[4\] u_cpu.rf_ram.memory\[113\]\[4\] u_cpu.rf_ram.memory\[114\]\[4\]
+ u_cpu.rf_ram.memory\[115\]\[4\] _01572_ _01573_ _01961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_20_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10418__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05086__A2 _01669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07050_ u_cpu.rf_ram.memory\[58\]\[4\] _03177_ _03182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06001_ _02463_ _02507_ _02508_ _02509_ _00072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_127_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09710__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06035__A1 _02402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10568__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06586__A2 u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07783__A1 _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07952_ u_cpu.rf_ram.memory\[120\]\[2\] _03693_ _03698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06903_ _02895_ _03089_ _03096_ _00387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09860__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09524__A2 _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07883_ u_cpu.rf_ram.memory\[92\]\[5\] _03652_ _03658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06338__A2 _02756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09622_ u_cpu.rf_ram.memory\[98\]\[1\] _04802_ _04804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06834_ _02768_ _02825_ _03058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09553_ _04628_ _04762_ _04765_ _01369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09288__A1 _04440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06765_ u_cpu.rf_ram.memory\[76\]\[1\] _03018_ _03020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05561__A3 _02139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08504_ _03896_ _04101_ _04106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05716_ u_cpu.cpu.mem_bytecnt\[1\] u_cpu.cpu.state.o_cnt\[2\] _02291_ _02292_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__07838__A2 _03626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09484_ _04636_ _04711_ _04718_ _01347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06696_ _02887_ _02978_ _02981_ _00295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08435_ u_cpu.rf_ram.memory\[114\]\[5\] _04041_ _04047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05647_ _01554_ _02224_ _01579_ _02225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_12_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06510__A2 _02861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08366_ _03899_ _03930_ _03988_ _03972_ _03989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05578_ _01617_ _02156_ _01600_ _02157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_109_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07317_ _03322_ _03325_ _03333_ _00564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10098__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09460__A1 _04630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08263__A2 _03885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08297_ u_arbiter.i_wb_cpu_rdt\[7\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[7\]
+ _02464_ _03925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06274__A1 _02685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07248_ u_cpu.rf_ram.memory\[140\]\[4\] _03287_ _03292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09212__A1 _04434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08015__A2 _03730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05872__I1 u_arbiter.i_wb_cpu_dbus_dat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07179_ _02657_ _03247_ _03253_ _00506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_65_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10190_ _00576_ io_in[4] u_cpu.rf_ram.memory\[70\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06577__A2 _02900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08318__A3 _03945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09515__A2 u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06329__A2 _02756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07829__A2 _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06501__A2 _02851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09733__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09451__A1 _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08254__A2 _03885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06265__A1 _02677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05068__A2 _01651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10526_ _00899_ io_in[4] u_cpu.rf_ram.memory\[116\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10710__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10457_ _00830_ io_in[4] u_cpu.rf_ram.memory\[117\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09883__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08557__A3 _03962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10388_ _00761_ io_in[4] u_cpu.rf_ram.memory\[37\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06568__A2 _02900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07765__A1 _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10860__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09506__A2 _04723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11009_ _01378_ io_in[4] u_cpu.rf_ram.memory\[25\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04880_ _01438_ _01467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_93_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08190__A1 u_arbiter.i_wb_cpu_rdt\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08317__I0 u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06740__A2 _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06550_ _02887_ _02883_ _02888_ _00242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06557__I _02656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05501_ _01638_ _02080_ _01482_ _02081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06481_ _02691_ _02840_ _02847_ _00214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09690__A1 _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05146__I3 u_cpu.rf_ram.memory\[139\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08220_ u_arbiter.i_wb_cpu_rdt\[21\] _03807_ _03829_ u_arbiter.i_wb_cpu_dbus_dat\[22\]
+ _03867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10240__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05432_ u_cpu.rf_ram.memory\[12\]\[5\] u_cpu.rf_ram.memory\[13\]\[5\] u_cpu.rf_ram.memory\[14\]\[5\]
+ u_cpu.rf_ram.memory\[15\]\[5\] _01530_ _01532_ _02012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_105_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08151_ u_arbiter.i_wb_cpu_dbus_dat\[2\] u_arbiter.i_wb_cpu_dbus_dat\[0\] u_arbiter.i_wb_cpu_dbus_dat\[1\]
+ _02915_ _03817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_05363_ _01505_ _01943_ _01579_ _01944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09442__A1 _04630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08245__A2 _03835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06256__A1 _02687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05059__A2 _01643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07102_ u_cpu.rf_ram.memory\[55\]\[3\] _03207_ _03211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05294_ u_cpu.rf_ram.memory\[116\]\[3\] u_cpu.rf_ram.memory\[117\]\[3\] u_cpu.rf_ram.memory\[118\]\[3\]
+ u_cpu.rf_ram.memory\[119\]\[3\] _01576_ _01577_ _01876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_107_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08082_ _03695_ _03770_ _03772_ _00891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10390__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07033_ _02652_ _03167_ _03172_ _00441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_127_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06008__A1 _02456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06559__A2 _02883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08984_ _02626_ _02766_ _04435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07935_ u_cpu.rf_ram.memory\[117\]\[4\] _03682_ _03687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07866_ _03637_ _03648_ _00799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04990__A1 _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08181__A1 u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09605_ _02681_ _04792_ _04794_ _01392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_95_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06817_ _03048_ _03049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_44_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07797_ u_cpu.cpu.state.o_cnt_r\[3\] u_cpu.cpu.state.o_cnt\[2\] _03604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_43_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06731__A2 _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09536_ u_cpu.rf_ram.memory\[27\]\[3\] _04752_ _04756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06748_ _02885_ _03008_ _03010_ _00318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09467_ u_cpu.rf_ram.memory\[87\]\[7\] _04701_ _04709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09756__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09681__A1 _04630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06679_ _02889_ _02967_ _02971_ _00288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08418_ _03969_ _04022_ _03958_ _04036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07800__B _02396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09398_ _04670_ _04671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_8_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10733__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08349_ _02909_ u_arbiter.i_wb_cpu_rdt\[14\] _03973_ _03974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09433__A1 _02870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08236__A2 _03808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06798__A2 _03037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10311_ _00697_ io_in[4] u_cpu.rf_ram.memory\[22\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10883__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10242_ _00628_ io_in[4] u_cpu.rf_ram.memory\[49\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07747__A1 _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10173_ _00559_ io_in[4] u_cpu.rf_ram.memory\[73\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05222__A2 _01804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10113__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06970__A2 _03137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05990__B _02456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06722__A2 _02988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10263__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05781__I0 u_arbiter.i_wb_cpu_dbus_dat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09672__A1 _02677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05289__A2 _01870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09424__A1 _04630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06238__A1 _02687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07986__A1 _03707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06789__A2 _03028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10509_ _00882_ io_in[4] u_cpu.rf_ram.memory\[122\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06410__A1 _02669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05981_ u_cpu.cpu.ctrl.o_ibus_adr\[9\] _02488_ _02456_ _02494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08538__I0 u_arbiter.i_wb_cpu_rdt\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06961__A2 _03127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07720_ u_cpu.rf_ram.memory\[124\]\[7\] _03553_ _03561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04932_ _01474_ _01479_ _01517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__10606__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08163__A1 _02915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07651_ _03522_ _03523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_04863_ _01441_ u_cpu.cpu.bne_or_bge _01442_ _01450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_53_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09779__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07910__A1 _03494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06713__A2 _02988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06602_ u_cpu.cpu.state.genblk1.misalign_trap_sync_r _02393_ _02926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05405__B _01471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07582_ u_cpu.rf_ram.memory\[130\]\[5\] _03475_ _03481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09321_ _04622_ _04624_ _04625_ _01277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10756__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06533_ _02687_ _02872_ _02877_ _00236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_90_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09663__A1 _04630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06477__A1 _02687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09252_ _04440_ _04583_ _04586_ _01247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06464_ _02693_ _02829_ _02837_ _00207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08203_ _03854_ _03855_ _00929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05415_ _01986_ _01995_ _01996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09183_ u_cpu.rf_ram.memory\[99\]\[4\] _04543_ _04548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09415__A1 _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06395_ _02683_ _02794_ _02797_ _00178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08134_ _02913_ _03801_ _03802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05346_ _01920_ _01922_ _01924_ _01926_ _01541_ _01927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_135_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08065_ u_cpu.rf_ram.memory\[122\]\[2\] _03760_ _03763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05277_ _01490_ _01849_ _01858_ _01859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_108_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07016_ u_cpu.rf_ram.memory\[19\]\[5\] _03157_ _03163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10136__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07729__A1 _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06401__A1 _02689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08967_ u_cpu.rf_ram.memory\[97\]\[0\] _04425_ _04426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06952__A2 _03127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10286__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07918_ _03504_ _03672_ _03677_ _00822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08898_ u_cpu.rf_ram.memory\[2\]\[3\] _04371_ _04375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_57_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07849_ u_cpu.rf_ram.memory\[90\]\[7\] _03626_ _03634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06704__A2 _02978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10860_ _01229_ io_in[4] u_cpu.rf_ram.memory\[105\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09519_ _01477_ _02294_ _04745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_25_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09654__A1 _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10791_ _01160_ io_in[4] u_cpu.rf_ram.memory\[28\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05140__A1 _01492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09406__A1 _04630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07968__A1 _03707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08361__B _03912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11061__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10225_ _00611_ io_in[4] u_cpu.rf_ram.memory\[39\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10629__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08393__A1 _04000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07196__A2 _03257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10156_ _00542_ io_in[4] u_cpu.rf_ram.memory\[13\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06943__A2 _03117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09921__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04954__A1 _01513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10087_ _00481_ io_in[4] u_cpu.rf_ram.memory\[54\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08145__A1 _03802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10779__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05054__S1 _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09645__A1 _04630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10989_ _01358_ io_in[4] u_cpu.cpu.genblk3.csr.o_new_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10009__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06835__I _03058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07120__A2 _03217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05200_ u_cpu.rf_ram.memory\[124\]\[2\] u_cpu.rf_ram.memory\[125\]\[2\] u_cpu.rf_ram.memory\[126\]\[2\]
+ u_cpu.rf_ram.memory\[127\]\[2\] _01496_ _01594_ _01783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_8_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06180_ _02606_ u_cpu.rf_ram_if.wdata1_r\[6\] _02659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__10159__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07959__A1 _03701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05131_ u_cpu.rf_ram.memory\[64\]\[1\] u_cpu.rf_ram.memory\[65\]\[1\] u_cpu.rf_ram.memory\[66\]\[1\]
+ u_cpu.rf_ram.memory\[67\]\[1\] _01522_ _01622_ _01715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_117_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05062_ _01637_ _01640_ _01644_ _01646_ _01466_ _01647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__06631__A1 _02897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09870_ _00264_ io_in[4] u_cpu.rf_ram.memory\[16\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08698__S _04257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07187__A2 _03257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08821_ _04331_ _01071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05198__A1 _01566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06934__A2 _03117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08752_ u_arbiter.i_wb_cpu_dbus_adr\[31\] _04290_ _02335_ _04291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05964_ u_cpu.cpu.ctrl.o_ibus_adr\[5\] _02476_ _02480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08136__A1 _03802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07703_ _03510_ _03543_ _03551_ _00732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_04915_ _01499_ _01500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08683_ u_cpu.rf_ram.memory\[31\]\[6\] _04247_ _04254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05895_ u_arbiter.i_wb_cpu_rdt\[18\] u_arbiter.i_wb_cpu_dbus_dat\[15\] _02431_ _02434_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08687__A2 _02392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06698__A1 _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07634_ u_cpu.rf_ram.memory\[128\]\[0\] _03513_ _03514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05370__A1 _01548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07565_ _03318_ _03465_ _03471_ _00674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09636__A1 _02717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08439__A2 _04041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04974__B _01558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09304_ _04438_ _04613_ _04615_ _01270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06516_ _02689_ _02861_ _02867_ _00229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07496_ u_cpu.rf_ram.memory\[135\]\[7\] _03425_ _03433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07111__A2 _03207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09235_ u_cpu.rf_ram.memory\[106\]\[3\] _04573_ _04577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06447_ _02825_ _02827_ _02828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09166_ _04444_ _04533_ _04538_ _01209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06870__A1 _02695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05673__A2 _02250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06378_ u_cpu.rf_ram.memory\[42\]\[3\] _02784_ _02788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11084__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08117_ u_cpu.rf_ram.memory\[33\]\[1\] _03790_ _03792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05329_ u_cpu.rf_ram.memory\[28\]\[4\] u_cpu.rf_ram.memory\[29\]\[4\] u_cpu.rf_ram.memory\[30\]\[4\]
+ u_cpu.rf_ram.memory\[31\]\[4\] _01497_ _01501_ _01910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09097_ u_arbiter.i_wb_cpu_rdt\[30\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[14\]
+ _04485_ _04500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08611__A2 u_arbiter.i_wb_cpu_rdt\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08048_ _03697_ _03750_ _03753_ _00876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09944__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08375__A1 _03974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07178__A2 _03247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10010_ _00404_ io_in[4] u_cpu.rf_ram.memory\[63\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08401__S _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05189__A1 _01490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09999_ _00393_ io_in[4] u_cpu.rf_ram.memory\[29\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06925__A2 _03100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10921__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08678__A2 _04247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10912_ _01281_ io_in[4] u_cpu.rf_ram.memory\[84\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05045__B _01481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06689__A1 _02695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07350__A2 _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10843_ _01212_ io_in[4] u_cpu.rf_ram.memory\[104\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09627__A1 _04630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05361__A1 _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10774_ _01143_ io_in[4] u_cpu.rf_ram.memory\[95\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07102__A2 _03207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10301__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05113__A1 _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06861__A1 _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05664__A2 _02241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08602__A2 _03986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10451__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08366__A1 _03899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07169__A2 _03247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08366__B2 _03972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10208_ _00594_ io_in[4] u_cpu.rf_ram.memory\[14\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06916__A2 _03100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10139_ _00525_ io_in[4] u_cpu.rf_ram.memory\[141\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05734__I _01442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08118__A1 _03695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08669__A2 _02870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05680_ _01473_ _02208_ _02257_ _00007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07341__A2 _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09618__A1 _02619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05352__A1 _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07350_ u_cpu.rf_ram.memory\[70\]\[6\] _03345_ _03352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09817__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06301_ u_cpu.rf_ram.memory\[1\]\[6\] _02733_ _02740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05104__A1 _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07281_ _03310_ _03308_ _03311_ _00550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09020_ _04444_ _04453_ _04458_ _01143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05655__A2 _02232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06852__A1 _02619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06232_ _02681_ _02697_ _02699_ _00113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06163_ _02611_ u_cpu.rf_ram_if.wdata0_r\[3\] _02644_ _02645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09967__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05114_ u_cpu.rf_ram.memory\[120\]\[1\] u_cpu.rf_ram.memory\[121\]\[1\] u_cpu.rf_ram.memory\[122\]\[1\]
+ u_cpu.rf_ram.memory\[123\]\[1\] _01598_ _01556_ _01698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_102_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05407__A2 _01987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06604__A1 _02912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06094_ _02305_ u_cpu.cpu.decode.opcode\[1\] _02584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10944__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09922_ _00316_ io_in[4] u_cpu.rf_ram.memory\[77\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05045_ _01512_ _01629_ _01481_ _01630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_113_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08357__A1 _03969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09853_ _00247_ io_in[4] u_cpu.rf_ram.memory\[50\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06907__A2 _02803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08804_ u_cpu.cpu.ctrl.o_ibus_adr\[10\] _04309_ _04311_ u_cpu.cpu.ctrl.o_ibus_adr\[11\]
+ _04322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_58_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09784_ _00178_ io_in[4] u_cpu.rf_ram.memory\[46\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__04918__A1 _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06996_ u_cpu.rf_ram.memory\[60\]\[4\] _03147_ _03152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07580__A2 _03475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08735_ _04280_ _01036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05947_ _02466_ _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_45_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05591__A1 _02160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05018__S1 _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08666_ _03705_ _04237_ _04244_ _01003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05878_ u_arbiter.i_wb_cpu_rdt\[10\] u_arbiter.i_wb_cpu_dbus_dat\[7\] _02418_ _02425_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_54_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07332__A2 _03335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10324__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07617_ _02646_ _03502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05343__A1 _01528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08597_ _03972_ _03985_ _04188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_26_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09609__A1 _02685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07548_ u_cpu.rf_ram.memory\[132\]\[6\] _03455_ _03462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07479_ _03322_ _03415_ _03423_ _00636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08832__A2 _04327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10474__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09218_ _04442_ _04563_ _04567_ _01232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06843__A1 _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10490_ _00863_ io_in[4] u_cpu.rf_ram.memory\[8\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09149_ u_cpu.rf_ram.memory\[103\]\[5\] _04523_ _04529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07399__A2 _03375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08596__A1 _03932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11111_ _00041_ io_in[0] u_arbiter.i_wb_cpu_rdt\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08348__A1 _02465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11042_ _01411_ io_in[4] u_cpu.rf_ram.memory\[100\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08899__A2 _04371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07020__A1 u_cpu.rf_ram.memory\[19\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05421__I2 u_cpu.rf_ram.memory\[22\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07323__A2 _03335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05334__A1 _01513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10826_ _01195_ io_in[4] u_cpu.rf_ram.memory\[102\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10817__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07087__A1 _03108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10757_ _01126_ io_in[4] u_cpu.rf_ram.memory\[97\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06834__A1 _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05193__S0 _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10688_ _01058_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08533__C _03910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10967__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08587__A1 _03924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05496__S1 _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07011__A1 _03104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06850_ u_cpu.rf_ram.memory\[67\]\[7\] _03059_ _03067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05801_ _02272_ _02371_ _02372_ _00016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07562__A2 _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10347__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06781_ u_cpu.rf_ram.memory\[75\]\[0\] _03028_ _03029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08520_ _04057_ _04119_ _04120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05732_ u_cpu.cpu.genblk3.csr.o_new_irq u_cpu.cpu.state.init_done _02307_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08511__A1 _03944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06117__A3 u_cpu.cpu.immdec.imm11_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07314__A2 _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08451_ _03925_ _03918_ _03988_ _03941_ _04060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_36_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05325__A1 _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05663_ u_cpu.rf_ram.memory\[72\]\[7\] u_cpu.rf_ram.memory\[73\]\[7\] u_cpu.rf_ram.memory\[74\]\[7\]
+ u_cpu.rf_ram.memory\[75\]\[7\] _01562_ _01563_ _02241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_51_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10497__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07402_ u_cpu.rf_ram.memory\[138\]\[5\] _03375_ _03381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05413__B _01482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08382_ _02285_ _03956_ _04003_ _00960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05594_ _01513_ _02171_ _02172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09067__A2 _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07333_ _03320_ _03335_ _03342_ _00571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_91_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06825__A1 _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07264_ u_cpu.rf_ram.memory\[13\]\[3\] _03297_ _03301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05184__S0 _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09003_ _02661_ _04448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06215_ u_cpu.rf_ram.memory\[21\]\[4\] _02679_ _02688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07195_ _02652_ _03257_ _03262_ _00513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__04931__S0 _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06146_ _02630_ _02631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06077_ u_cpu.cpu.ctrl.o_ibus_adr\[28\] u_cpu.cpu.ctrl.o_ibus_adr\[27\] _02562_ _02571_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__05487__S1 _01563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11122__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05028_ u_cpu.rf_ram.memory\[88\]\[0\] u_cpu.rf_ram.memory\[89\]\[0\] u_cpu.rf_ram.memory\[90\]\[0\]
+ u_cpu.rf_ram.memory\[91\]\[0\] _01598_ _01577_ _01613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_99_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09905_ _00299_ io_in[4] u_cpu.rf_ram.memory\[129\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09836_ _00230_ io_in[4] u_cpu.rf_ram.memory\[48\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08750__A1 u_cpu.cpu.bufreg.i_sh_signed vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09767_ _00161_ io_in[4] u_cpu.rf_ram.memory\[78\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06979_ _03108_ _03137_ _03142_ _00417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08718_ u_arbiter.i_wb_cpu_dbus_adr\[16\] u_arbiter.i_wb_cpu_dbus_adr\[17\] _04257_
+ _04272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_26_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09698_ _04845_ _01434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08502__A1 u_cpu.cpu.immdec.imm30_25\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07305__A2 _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05316__A1 _01492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08649_ u_cpu.cpu.genblk3.csr.mie_mtie u_cpu.cpu.genblk3.csr.mstatus_mie u_cpu.cpu.genblk3.csr.i_mtip
+ _04234_ _04235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_55_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09058__A2 _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10611_ _00984_ io_in[4] u_cpu.cpu.immdec.imm30_25\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07069__A1 _03108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08634__B _03969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10542_ _00915_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06816__A1 _02717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05175__S0 _01551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06292__A2 _02733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10473_ _00846_ io_in[4] u_cpu.rf_ram.memory\[118\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09230__A2 _04573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07241__A1 _03098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05993__B _02461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05478__S1 _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07792__A2 _03593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11025_ _01394_ io_in[4] u_cpu.rf_ram.memory\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07544__A2 _03455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05555__A1 _01566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04989__S0 _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05650__S1 _01563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09297__A2 _04603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05858__A2 _02403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05233__B _01534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10809_ _01178_ io_in[4] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06807__A1 _02647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05166__S0 _01523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07480__A1 _02743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11145__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06000_ _02402_ u_scanchain_local.module_data_in\[50\] _02478_ u_arbiter.i_wb_cpu_dbus_adr\[13\]
+ _02509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__05491__B1 _02068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09221__A2 _04563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08980__A1 _03705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07783__A2 _03593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07951_ _02641_ _03697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05794__A1 _01460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06902_ u_cpu.rf_ram.memory\[64\]\[6\] _03089_ _03096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07882_ _03504_ _03652_ _03657_ _00806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09621_ _04622_ _04802_ _04803_ _01399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06833_ _02897_ _03049_ _03057_ _00356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05546__A1 _01548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09552_ u_cpu.rf_ram.memory\[26\]\[2\] _04762_ _04765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06764_ _02881_ _03018_ _03019_ _00325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09288__A2 _04603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08503_ _04098_ _04103_ _04105_ _00979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05715_ u_cpu.cpu.mem_bytecnt\[0\] _02291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07299__A1 _03322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09483_ u_cpu.rf_ram.memory\[88\]\[6\] _04711_ _04718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06695_ u_cpu.rf_ram.memory\[129\]\[2\] _02978_ _02981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08434_ _03701_ _04041_ _04046_ _00969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05646_ u_cpu.rf_ram.memory\[116\]\[7\] u_cpu.rf_ram.memory\[117\]\[7\] u_cpu.rf_ram.memory\[118\]\[7\]
+ u_cpu.rf_ram.memory\[119\]\[7\] _01576_ _01577_ _02224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_93_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08365_ _03974_ _03908_ _03988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05577_ u_cpu.rf_ram.memory\[76\]\[6\] u_cpu.rf_ram.memory\[77\]\[6\] u_cpu.rf_ram.memory\[78\]\[6\]
+ u_cpu.rf_ram.memory\[79\]\[6\] _01529_ _01500_ _02156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07316_ u_cpu.rf_ram.memory\[73\]\[7\] _03325_ _03333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05157__S0 _01497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08296_ u_arbiter.i_wb_cpu_rdt\[9\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[9\]
+ _02464_ _03924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09460__A2 _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06274__A2 _02719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07247_ _03106_ _03287_ _03291_ _00536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07471__A1 _03314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07178_ u_cpu.rf_ram.memory\[9\]\[5\] _03247_ _03253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09212__A2 _04563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10512__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07223__A1 _03098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06129_ _02609_ _02613_ _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_65_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07774__A2 _03583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08318__A4 _03899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09515__A3 _02291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10662__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07526__A2 _03445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09819_ _00213_ io_in[4] u_cpu.rf_ram.memory\[41\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05537__A1 _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09279__A2 _04593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11018__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10042__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05148__S0 _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09451__A2 _02743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06265__A2 _02717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10525_ _00898_ io_in[4] u_cpu.rf_ram.memory\[116\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07462__A1 _02954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10456_ _00829_ io_in[4] u_cpu.rf_ram.memory\[117\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09203__A2 _04553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10192__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10387_ _00760_ io_in[4] u_cpu.rf_ram.memory\[37\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08962__A1 _03956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07765__A2 _03583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04911__I _01495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05320__S0 _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11008_ _01377_ io_in[4] u_cpu.rf_ram.memory\[25\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05528__A1 _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08539__B _03922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08190__A2 _03822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08317__I1 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05500_ u_cpu.rf_ram.memory\[132\]\[5\] u_cpu.rf_ram.memory\[133\]\[5\] u_cpu.rf_ram.memory\[134\]\[5\]
+ u_cpu.rf_ram.memory\[135\]\[5\] _01641_ _01642_ _02080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_34_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06480_ u_cpu.rf_ram.memory\[41\]\[6\] _02840_ _02847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09690__A2 _03611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05431_ _01528_ _02010_ _02011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08150_ u_arbiter.i_wb_cpu_dbus_dat\[3\] _02915_ _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05362_ u_cpu.rf_ram.memory\[48\]\[4\] u_cpu.rf_ram.memory\[49\]\[4\] u_cpu.rf_ram.memory\[50\]\[4\]
+ u_cpu.rf_ram.memory\[51\]\[4\] _01576_ _01577_ _01943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09442__A2 _04691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10535__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07101_ _03104_ _03207_ _03210_ _00471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08081_ u_cpu.rf_ram.memory\[115\]\[1\] _03770_ _03772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06256__A2 _02707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07453__A1 _03314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05293_ _01602_ _01874_ _01875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07032_ u_cpu.rf_ram.memory\[5\]\[4\] _03167_ _03172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_127_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07205__A1 _03098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10685__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08953__A1 u_cpu.cpu.immdec.imm11_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07756__A2 _03573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05767__A1 _02305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05311__S0 _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08983_ _02631_ _04434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07934_ _03502_ _03682_ _03686_ _00829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05138__B _01481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07508__A2 _03435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07865_ _02265_ _03647_ _00773_ _02305_ _03648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__05519__A1 _01528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08449__B _03975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08181__A2 _03822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09604_ u_cpu.rf_ram.memory\[0\]\[1\] _04792_ _04794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_28_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06816_ _02717_ _02768_ _03048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07796_ _03603_ _00773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_3_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09535_ _04628_ _04752_ _04755_ _01361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06747_ u_cpu.rf_ram.memory\[74\]\[1\] _03008_ _03010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09130__A1 _04444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10065__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09466_ _04636_ _04701_ _04708_ _01339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06678_ u_cpu.rf_ram.memory\[119\]\[3\] _02967_ _02971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05378__S0 _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09681__A2 _04832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06495__A2 _02851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08417_ _03986_ _04034_ _04035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05629_ _01489_ _02197_ _02206_ _02207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_09397_ _02766_ _04349_ _04670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08348_ _02465_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[14\] _03973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_138_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09433__A2 _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06247__A2 _02707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07444__A1 _02695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08279_ _02465_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\] _03907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_138_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10310_ _00696_ io_in[4] u_cpu.rf_ram.memory\[22\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07995__A2 _03720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10241_ _00627_ io_in[4] u_cpu.rf_ram.memory\[49\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05058__I0 u_cpu.rf_ram.memory\[128\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08944__A1 _03945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07747__A2 _03573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10172_ _00558_ io_in[4] u_cpu.rf_ram.memory\[73\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05302__S0 _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05048__B _01471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10408__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05930__A1 _02403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05781__I1 u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05369__S0 _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09672__A2 _02743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10558__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07683__A1 _03508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04906__I _01467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09850__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09424__A2 _04681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07435__A1 _03314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06238__A2 _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07986__A2 _03710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10508_ _00881_ io_in[4] u_cpu.rf_ram.memory\[112\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05997__A1 _02389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09188__A1 _04448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10439_ _00812_ io_in[4] u_cpu.rf_ram.memory\[35\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07738__A2 _03563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08935__B2 _03910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05749__A1 _02322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06410__A2 _02805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05980_ _02492_ _02486_ _02487_ _02493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_111_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08538__I1 u_arbiter.i_wb_cpu_rdt\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04931_ u_cpu.rf_ram.memory\[16\]\[0\] u_cpu.rf_ram.memory\[17\]\[0\] u_cpu.rf_ram.memory\[18\]\[0\]
+ u_cpu.rf_ram.memory\[19\]\[0\] _01508_ _01509_ _01516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_111_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10088__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09360__A1 _04638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07650_ _02870_ _02965_ _03522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04862_ _01448_ u_cpu.cpu.decode.op26 u_cpu.cpu.decode.co_ebreak _01449_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_65_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06174__A1 _02606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06601_ _02313_ _02923_ _02924_ _02925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07910__A2 _03672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07581_ _03316_ _03475_ _03480_ _00681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09112__A1 _04444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09320_ u_cpu.rf_ram.memory\[84\]\[0\] _04624_ _04625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06532_ u_cpu.rf_ram.memory\[47\]\[4\] _02872_ _02877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09663__A2 _04822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09251_ u_cpu.rf_ram.memory\[107\]\[2\] _04583_ _04586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06477__A2 _02840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06463_ u_cpu.rf_ram.memory\[51\]\[7\] _02829_ _02837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08202_ u_arbiter.i_wb_cpu_rdt\[15\] _03822_ _03833_ u_arbiter.i_wb_cpu_dbus_dat\[16\]
+ _03855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_21_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05414_ _01988_ _01990_ _01992_ _01994_ _01466_ _01995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_09182_ _04442_ _04543_ _04547_ _01216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06394_ u_cpu.rf_ram.memory\[46\]\[2\] _02794_ _02797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09415__A2 _03037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08133_ _02259_ _03799_ _03800_ _03801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_105_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05345_ _01513_ _01925_ _01482_ _01926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07426__A1 _02838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06229__A2 _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07977__A2 _03710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08064_ _03695_ _03760_ _03762_ _00883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05276_ _01851_ _01853_ _01855_ _01857_ _01581_ _01858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__05532__S0 _01496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07015_ _03108_ _03157_ _03162_ _00433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07729__A2 _03563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08926__A1 _02392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06401__A2 _02794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08966_ _04424_ _04425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_64_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07917_ u_cpu.rf_ram.memory\[34\]\[4\] _03672_ _03677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08897_ _02642_ _04371_ _04374_ _01104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09723__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07848_ _03508_ _03626_ _03633_ _00795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05599__S0 _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07901__A2 _03662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05315__C _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10700__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07779_ _03494_ _03593_ _03594_ _00765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09518_ _04741_ _04743_ _04744_ _01355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10790_ _01159_ io_in[4] u_cpu.rf_ram.memory\[28\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09873__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09654__A2 _02838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07665__A1 _03508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06468__A2 _02840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09449_ u_cpu.rf_ram.memory\[111\]\[7\] _04691_ _04699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10850__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09406__A2 _04671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07417__A1 _03314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07968__A2 _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08090__A1 _03703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05523__S0 _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06640__A2 _02945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05294__I3 u_cpu.rf_ram.memory\[119\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08917__A1 _03699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10224_ _00610_ io_in[4] u_cpu.rf_ram.memory\[39\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10155_ _00541_ io_in[4] u_cpu.rf_ram.memory\[13\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10230__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10086_ _00480_ io_in[4] u_cpu.rf_ram.memory\[54\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09342__A1 _04638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06156__A1 _02606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10380__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09645__A2 _04812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10988_ _01357_ io_in[4] u_cpu.cpu.ctrl.i_iscomp vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06459__A2 _02829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07408__A1 _02743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07959__A2 _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05130_ _01707_ _01709_ _01711_ _01713_ _01486_ _01714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_116_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05514__S0 _01523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06092__B1 _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05061_ _01638_ _01645_ _01482_ _01646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06631__A2 _02935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06072__B _02397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08908__A1 _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08384__A2 _04004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09746__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09581__A1 _04638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08820_ u_cpu.cpu.ctrl.o_ibus_adr\[17\] _04327_ _04329_ u_cpu.cpu.ctrl.o_ibus_adr\[18\]
+ _04331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06395__A1 _02683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05963_ _02463_ _02477_ _02479_ _00063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08751_ _04288_ _04289_ _04290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10723__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09333__A1 _04632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07702_ u_cpu.rf_ram.memory\[125\]\[7\] _03543_ _03551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04914_ _01498_ _01499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08682_ _03703_ _04247_ _04253_ _01010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05894_ _02433_ _00038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09896__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06698__A2 _02978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07633_ _03512_ _03513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_54_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07564_ u_cpu.rf_ram.memory\[131\]\[5\] _03465_ _03471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10873__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09636__A2 _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06515_ u_cpu.rf_ram.memory\[48\]\[5\] _02861_ _02867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09303_ u_cpu.rf_ram.memory\[69\]\[1\] _04613_ _04615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07647__A1 _03508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07495_ _03320_ _03425_ _03432_ _00643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08844__B1 _04329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09234_ _04440_ _04573_ _04576_ _01239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06446_ _02826_ _02827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10103__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09165_ u_cpu.rf_ram.memory\[104\]\[4\] _04533_ _04538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06870__A2 _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06377_ _02683_ _02784_ _02787_ _00170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08116_ _03691_ _03790_ _03791_ _00906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__04881__A1 u_cpu.cpu.immdec.imm19_12_20\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05328_ _01473_ _01860_ _01909_ _00003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_134_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08072__A1 _03703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09096_ _04499_ _01178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05505__S0 _01497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08047_ u_cpu.rf_ram.memory\[112\]\[2\] _03750_ _03753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06622__A2 _02935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05259_ u_cpu.rf_ram.memory\[36\]\[3\] u_cpu.rf_ram.memory\[37\]\[3\] u_cpu.rf_ram.memory\[38\]\[3\]
+ u_cpu.rf_ram.memory\[39\]\[3\] _01544_ _01545_ _01841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10253__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08375__A2 _03947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05189__A2 _01762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09998_ _00392_ io_in[4] u_cpu.rf_ram.memory\[29\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08949_ _02728_ _04390_ _04411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09324__A1 _04626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08127__A2 _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06138__A1 _02621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10911_ _01280_ io_in[4] u_cpu.rf_ram.memory\[84\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07886__A1 _03508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06689__A2 _02976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10842_ _01211_ io_in[4] u_cpu.rf_ram.memory\[104\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05361__A2 _01941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09627__A2 _04802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08356__C _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10773_ _01142_ io_in[4] u_cpu.rf_ram.memory\[95\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05061__B _01482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05113__A2 _01696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06310__A1 _02632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06861__A2 _03069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04872__A1 u_cpu.cpu.decode.op21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09769__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07810__A1 _02396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10746__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09563__A1 _04638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10207_ _00593_ io_in[4] u_cpu.rf_ram.memory\[14\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06377__A1 _02683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10138_ _00524_ io_in[4] u_cpu.rf_ram.memory\[142\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08118__A2 _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10069_ _00463_ io_in[4] u_cpu.rf_ram.memory\[56\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10896__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09618__A2 _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05750__I u_cpu.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05352__A2 _01932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10126__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08826__B1 _04329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06300_ _02657_ _02733_ _02739_ _00141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07280_ u_cpu.rf_ram.memory\[72\]\[1\] _03308_ _03311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06231_ u_cpu.rf_ram.memory\[81\]\[1\] _02697_ _02699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06852__A2 _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10276__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04863__A1 _01441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08054__A1 _03703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06162_ _02606_ u_cpu.rf_ram_if.wdata1_r\[3\] _02644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_117_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05113_ _01543_ _01696_ _01697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06604__A2 _02927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06093_ _02463_ _02582_ _02583_ _00091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07801__A1 _02291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05044_ u_cpu.rf_ram.memory\[76\]\[0\] u_cpu.rf_ram.memory\[77\]\[0\] u_cpu.rf_ram.memory\[78\]\[0\]
+ u_cpu.rf_ram.memory\[79\]\[0\] _01529_ _01500_ _01629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09921_ _00315_ io_in[4] u_cpu.rf_ram.memory\[77\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09852_ _00246_ io_in[4] u_cpu.rf_ram.memory\[50\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06368__A1 u_cpu.cpu.immdec.imm11_7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08803_ _04321_ _01063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_86_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09783_ _00177_ io_in[4] u_cpu.rf_ram.memory\[46\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__04918__A2 _01502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06995_ _03106_ _03147_ _03151_ _00424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08109__A2 _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09306__A1 _04440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08734_ u_arbiter.i_wb_cpu_dbus_adr\[24\] u_arbiter.i_wb_cpu_dbus_adr\[25\] _02335_
+ _04280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_100_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05946_ _02465_ _02466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05591__A2 _02169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05877_ _02424_ _00029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08665_ u_cpu.rf_ram.memory\[32\]\[6\] _04237_ _04244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08457__B _03966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04985__B _01480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07616_ _03500_ _03496_ _03501_ _00695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08596_ _03932_ _03906_ _04031_ _04051_ _04187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__05343__A2 _01923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09609__A2 _04792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11051__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07547_ _03318_ _03455_ _03461_ _00666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10619__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08293__A1 _02464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07478_ u_cpu.rf_ram.memory\[136\]\[7\] _03415_ _03423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07096__A2 _03207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09217_ u_cpu.rf_ram.memory\[105\]\[3\] _04563_ _04567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06843__A2 _03059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06429_ _02669_ _02816_ _02817_ _00192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09911__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09148_ _04444_ _04523_ _04528_ _01201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09093__I0 u_arbiter.i_wb_cpu_rdt\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10769__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08596__A2 _03906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09079_ u_arbiter.i_wb_cpu_rdt\[21\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[5\]
+ _04485_ _04491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11110_ _00040_ io_in[0] u_arbiter.i_wb_cpu_rdt\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08412__S _02466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11041_ _01410_ io_in[4] u_cpu.rf_ram.memory\[100\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09545__A1 _04638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06359__A1 _02687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05835__I io_in[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07020__A2 _03157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05031__A1 _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10149__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06531__A1 _02685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10825_ _01194_ io_in[4] u_cpu.rf_ram.memory\[102\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08808__B1 _04311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10299__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08284__A1 _03904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07087__A2 _03197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10756_ _01125_ io_in[4] u_cpu.rf_ram.memory\[97\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06834__A2 _02825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10687_ _01057_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05193__S1 _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05893__I0 u_arbiter.i_wb_cpu_rdt\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08036__A1 _02657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04914__I _01498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08587__A2 _04052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07011__A2 _03157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05800_ _02272_ u_cpu.rf_ram_if.rdata1\[2\] _02372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06780_ _03027_ _03028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06770__A1 _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07960__I _02656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05731_ u_cpu.cpu.bufreg.lsb\[0\] _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11074__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08511__A2 _03975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05662_ _01617_ _02239_ _01607_ _02240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08450_ _03980_ _03929_ _04058_ _04059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_91_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06522__A1 _02782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07401_ _03316_ _03375_ _03380_ _00601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_63_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08381_ _03965_ _03972_ _03994_ _04002_ _03955_ _04003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_05593_ u_cpu.rf_ram.memory\[28\]\[7\] u_cpu.rf_ram.memory\[29\]\[7\] u_cpu.rf_ram.memory\[30\]\[7\]
+ u_cpu.rf_ram.memory\[31\]\[7\] _01497_ _01501_ _02171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09934__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07332_ u_cpu.rf_ram.memory\[71\]\[6\] _03335_ _03342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08275__A1 _02465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07078__A2 _03197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07263_ _02642_ _03297_ _03300_ _00543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10911__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06825__A2 _03049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05184__S1 _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09002_ _04446_ _04436_ _04447_ _01136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05884__I0 u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06214_ _02651_ _02687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09075__I0 u_arbiter.i_wb_cpu_rdt\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07194_ u_cpu.rf_ram.memory\[15\]\[4\] _03257_ _03262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04931__S1 _01509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06145_ u_cpu.rf_ram_if.wdata0_r\[0\] _02611_ _02629_ _02630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_117_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06589__A1 _01444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06076_ u_cpu.cpu.ctrl.o_ibus_adr\[27\] _02562_ u_cpu.cpu.ctrl.o_ibus_adr\[28\] _02570_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07250__A2 _03287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09527__A1 _02395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05027_ _01464_ _01611_ _01612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09904_ _00298_ io_in[4] u_cpu.rf_ram.memory\[129\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07002__A2 _03147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09835_ _00229_ io_in[4] u_cpu.rf_ram.memory\[48\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08750__A2 u_arbiter.i_wb_cpu_dbus_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09766_ _00160_ io_in[4] u_cpu.rf_ram.memory\[78\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_101_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06761__A1 _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06978_ u_cpu.rf_ram.memory\[61\]\[4\] _03137_ _03142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08717_ _04271_ _01027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05929_ u_arbiter.i_wb_cpu_dbus_dat\[31\] _02452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09697_ _02396_ u_cpu.rf_ram_if.rreq_r _04845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_54_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08648_ _02263_ _02598_ _04234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10441__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08579_ u_cpu.cpu.csr_imm _03897_ _04164_ _04172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10610_ _00983_ io_in[4] u_cpu.cpu.immdec.imm30_25\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08266__A1 _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07069__A2 _03187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10591__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10541_ _00914_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06816__A2 _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05175__S1 _01524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08018__A1 _02657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10472_ _00845_ io_in[4] u_cpu.rf_ram.memory\[118\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07241__A2 _03287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09807__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11024_ _01393_ io_in[4] u_cpu.rf_ram.memory\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11097__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04989__S1 _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06752__A1 _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09957__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10934__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08257__A1 _03699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10808_ _01177_ io_in[4] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08317__S _02466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06807__A2 _03039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10739_ _01108_ io_in[4] u_cpu.rf_ram.memory\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05166__S1 _01525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05866__I0 u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07480__A2 _02976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07232__A2 _03277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10314__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08980__A2 _04425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07950_ _03695_ _03693_ _03696_ _00835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06991__A1 _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06901_ _02893_ _03089_ _03095_ _00386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07881_ u_cpu.rf_ram.memory\[92\]\[4\] _03652_ _03657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08193__B1 _03833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09620_ u_cpu.rf_ram.memory\[98\]\[0\] _04802_ _04803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06832_ u_cpu.rf_ram.memory\[68\]\[7\] _03049_ _03057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10464__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06743__A1 _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09551_ _04626_ _04762_ _04764_ _01368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06763_ u_cpu.rf_ram.memory\[76\]\[0\] _03018_ _03019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08502_ u_cpu.cpu.immdec.imm30_25\[0\] _04104_ _04105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05424__B _01519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05714_ u_cpu.cpu.decode.op22 _02290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09482_ _04634_ _04711_ _04717_ _01346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06694_ _02885_ _02978_ _02980_ _00294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07299__A2 _03308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08433_ u_cpu.rf_ram.memory\[114\]\[4\] _04041_ _04046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05645_ _01505_ _02222_ _02223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08248__A1 _02695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05576_ _01621_ _02154_ _02155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08364_ _03940_ _03941_ _03971_ _03987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08454__C _03938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07315_ _03320_ _03325_ _03332_ _00563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08295_ u_arbiter.i_wb_cpu_rdt\[10\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[10\]
+ _02464_ _03923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__05157__S1 _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07246_ u_cpu.rf_ram.memory\[140\]\[3\] _03287_ _03291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07471__A2 _03415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07177_ _02652_ _03247_ _03252_ _00505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_117_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06128_ _01460_ _02610_ _02612_ _02613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08420__A1 _04031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07223__A2 _03277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08971__A2 _04425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06059_ u_arbiter.i_wb_cpu_dbus_adr\[24\] _02397_ _02554_ _02556_ _02402_ _02557_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_120_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10807__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09515__A4 _02290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08184__B1 _03833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09818_ _00212_ io_in[4] u_cpu.rf_ram.memory\[41\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06734__A1 _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05537__A2 _02115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09749_ _00143_ io_in[4] u_cpu.rf_ram.memory\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10957__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08487__A1 _03966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08239__A1 u_arbiter.i_wb_cpu_dbus_dat\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05148__S1 _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10524_ _00897_ io_in[4] u_cpu.rf_ram.memory\[115\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07462__A2 _02976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10337__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05473__A1 _01490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10455_ _00828_ io_in[4] u_cpu.rf_ram.memory\[117\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08380__B _03969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07214__A2 _03267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10386_ _00759_ io_in[4] u_cpu.rf_ram.memory\[37\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08962__A2 _03922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10487__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05320__S1 _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06973__A1 _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08175__B1 _03833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11007_ _01376_ io_in[4] u_cpu.rf_ram.memory\[25\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06725__A1 _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05528__A2 _02106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05244__B _01481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08478__A1 _03912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06059__C _02402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05430_ u_cpu.rf_ram.memory\[8\]\[5\] u_cpu.rf_ram.memory\[9\]\[5\] u_cpu.rf_ram.memory\[10\]\[5\]
+ u_cpu.rf_ram.memory\[11\]\[5\] _01523_ _01525_ _02010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__11112__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05361_ _01571_ _01941_ _01942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07100_ u_cpu.rf_ram.memory\[55\]\[2\] _03207_ _03210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08080_ _03691_ _03770_ _03771_ _00890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05292_ u_cpu.rf_ram.memory\[112\]\[3\] u_cpu.rf_ram.memory\[113\]\[3\] u_cpu.rf_ram.memory\[114\]\[3\]
+ u_cpu.rf_ram.memory\[115\]\[3\] _01572_ _01545_ _01874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_9_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07453__A2 _03405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07031_ _02647_ _03167_ _03171_ _00440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08402__A1 _03944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07205__A2 _03267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08982_ _03707_ _04425_ _04433_ _01130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05311__S1 _01622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07933_ u_cpu.rf_ram.memory\[117\]\[3\] _03682_ _03686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07864_ _02286_ _03646_ _03647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_56_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06716__A1 _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09603_ _02669_ _04792_ _04793_ _01391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_95_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08449__C _03972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06815_ _02667_ _03039_ _03047_ _00348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_3_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07795_ _02395_ _03602_ _03603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09534_ u_cpu.rf_ram.memory\[27\]\[2\] _04752_ _04755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06746_ _02881_ _03008_ _03009_ _00317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08469__B2 _04039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09130__A2 _04513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09465_ u_cpu.rf_ram.memory\[87\]\[6\] _04701_ _04708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06677_ _02887_ _02967_ _02970_ _00287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_19_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07141__A1 _03108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05378__S1 _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08416_ _03974_ _04033_ _04024_ _03915_ _04034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_58_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05628_ _02199_ _02201_ _02203_ _02205_ _01485_ _02206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_09396_ _04638_ _04661_ _04669_ _01308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07692__A2 _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08347_ u_arbiter.i_wb_cpu_rdt\[13\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[13\]
+ _02466_ _03972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05559_ _01554_ _02137_ _01607_ _02138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05601__C _01486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08278_ _03905_ _03906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08641__A1 u_cpu.cpu.immdec.imm19_12_20\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07444__A2 _02827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07229_ _03106_ _03277_ _03281_ _00528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09197__A2 _04553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10240_ _00626_ io_in[4] u_cpu.rf_ram.memory\[49\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05207__A1 _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08944__A2 _03988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10171_ _00557_ io_in[4] u_cpu.rf_ram.memory\[73\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06955__A1 _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05302__S1 _01594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06707__A1 _02849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11135__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05781__I2 u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09121__A2 _04513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05369__S1 _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07683__A2 _03533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05694__A1 _02263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08632__A1 _04165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07435__A2 _03395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10507_ _00880_ io_in[4] u_cpu.rf_ram.memory\[112\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09188__A2 _04543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04922__I _01494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10438_ _00811_ io_in[4] u_cpu.rf_ram.memory\[35\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07199__A1 _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10369_ _00742_ io_in[4] u_cpu.rf_ram.memory\[123\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04930_ _01513_ _01514_ _01515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09360__A2 _04641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04861_ u_cpu.cpu.decode.op21 _01448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_93_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07371__A1 _03322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06600_ u_arbiter.i_wb_cpu_ack _02397_ _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07580_ u_cpu.rf_ram.memory\[130\]\[4\] _03475_ _03480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09112__A2 _04503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06531_ _02685_ _02872_ _02876_ _00235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10502__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07123__A1 _03108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09250_ _04438_ _04583_ _04585_ _01246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06584__I _02464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06462_ _02691_ _02829_ _02836_ _00206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08871__A1 _03707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07674__A2 _03533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08201_ u_arbiter.i_wb_cpu_dbus_dat\[15\] _03835_ _03854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05685__A1 u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05413_ _01638_ _01993_ _01482_ _01994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09181_ u_cpu.rf_ram.memory\[99\]\[3\] _04543_ _04547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06393_ _02681_ _02794_ _02796_ _00177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10652__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08132_ u_cpu.cpu.mem_bytecnt\[1\] _02355_ _03800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05344_ u_cpu.rf_ram.memory\[12\]\[4\] u_cpu.rf_ram.memory\[13\]\[4\] u_cpu.rf_ram.memory\[14\]\[4\]
+ u_cpu.rf_ram.memory\[15\]\[4\] _01530_ _01532_ _01925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08623__A1 _03923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07426__A2 _02976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08063_ u_cpu.rf_ram.memory\[122\]\[1\] _03760_ _03762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05275_ _01505_ _01856_ _01579_ _01857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05532__S1 _01594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09179__A2 _04543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07014_ u_cpu.rf_ram.memory\[19\]\[4\] _03157_ _03162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11008__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05149__B _01534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08926__A2 _02604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06937__A1 _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08965_ _02695_ _04349_ _04424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07916_ _03502_ _03672_ _03676_ _00821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10032__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08896_ u_cpu.rf_ram.memory\[2\]\[2\] _04371_ _04374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09351__A2 _04641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07847_ u_cpu.rf_ram.memory\[90\]\[6\] _03626_ _03633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05599__S1 _01509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07778_ u_cpu.rf_ram.memory\[36\]\[0\] _03593_ _03594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09071__S _04485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10182__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09103__A2 _04503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09517_ _02301_ _04743_ _02396_ _04744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06729_ u_cpu.rf_ram.memory\[77\]\[1\] _02998_ _03000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09448_ _04636_ _04691_ _04698_ _01331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07665__A2 _03523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09379_ _02626_ _02675_ _04660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05140__A3 _01723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07417__A2 _03385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08090__A2 _03770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05523__S1 _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08917__A2 _04381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10223_ _00609_ io_in[4] u_cpu.rf_ram.memory\[39\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06928__A1 _03112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09590__A2 _04782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10154_ _00540_ io_in[4] u_cpu.rf_ram.memory\[140\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05600__A1 _01506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10085_ _00479_ io_in[4] u_cpu.rf_ram.memory\[54\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09342__A2 _04624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10525__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07353__A1 _03322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10987_ _01356_ io_in[4] u_cpu.cpu.genblk3.csr.mstatus_mie vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07105__A1 _03108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10675__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07656__A2 _03523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08853__A1 u_cpu.cpu.immdec.imm11_7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07408__A2 _02782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__04890__A2 _01443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08081__A2 _03770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05514__S1 _01525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06092__A1 _02402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05060_ u_cpu.rf_ram.memory\[132\]\[0\] u_cpu.rf_ram.memory\[133\]\[0\] u_cpu.rf_ram.memory\[134\]\[0\]
+ u_cpu.rf_ram.memory\[135\]\[0\] _01641_ _01642_ _01645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_99_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06092__B2 u_arbiter.i_wb_cpu_dbus_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08369__B1 _03985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08908__A2 _02803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09030__A1 _04434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10055__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06919__A1 _03106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07963__I _02661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09581__A2 _04772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06395__A2 _02794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08750_ u_cpu.cpu.bufreg.i_sh_signed u_arbiter.i_wb_cpu_dbus_adr\[31\] _02598_ _04289_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05962_ _02403_ u_scanchain_local.module_data_in\[42\] _02478_ u_arbiter.i_wb_cpu_dbus_adr\[5\]
+ _02479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07701_ _03508_ _03543_ _03550_ _00731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09333__A2 _04624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04913_ u_cpu.raddr\[1\] _01498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08681_ u_cpu.rf_ram.memory\[31\]\[5\] _04247_ _04253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05893_ u_arbiter.i_wb_cpu_rdt\[17\] u_arbiter.i_wb_cpu_dbus_dat\[14\] _02431_ _02433_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_65_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07632_ _02754_ _02976_ _03512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07895__A2 _03662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05450__S0 _01576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07563_ _03316_ _03465_ _03470_ _00673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09302_ _04434_ _04613_ _04614_ _01269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06514_ _02687_ _02861_ _02866_ _00228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07494_ u_cpu.rf_ram.memory\[135\]\[6\] _03425_ _03432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07647__A2 _03513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05202__S0 _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09233_ u_cpu.rf_ram.memory\[106\]\[2\] _04573_ _04576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06445_ _02728_ u_cpu.cpu.immdec.imm11_7\[4\] _02622_ _02729_ _02826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_10_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09164_ _04442_ _04533_ _04537_ _01208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06376_ u_cpu.rf_ram.memory\[42\]\[2\] _02784_ _02787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08115_ u_cpu.rf_ram.memory\[33\]\[0\] _03790_ _03791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__04881__A2 _01467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05327_ _01899_ _01908_ _01909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08072__A2 _03760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09095_ u_arbiter.i_wb_cpu_rdt\[29\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[13\]
+ _04485_ _04499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__05505__S1 _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06083__A1 _02463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08046_ _03695_ _03750_ _03752_ _00875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05258_ _01833_ _01835_ _01837_ _01839_ _01541_ _01840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__05830__A1 io_in[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05189_ _01490_ _01762_ _01771_ _01772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09572__A2 _04772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09997_ _00391_ io_in[4] u_cpu.rf_ram.memory\[29\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10548__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05189__A3 _01771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07583__A1 _03318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06386__A2 _02784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08948_ _03896_ _04407_ _04409_ _04410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_48_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09840__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09324__A2 _04624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05326__C _01466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08879_ _02642_ _04361_ _04364_ _01096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_57_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06138__A2 _02622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07335__A1 _03322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10910_ _01279_ io_in[4] u_cpu.rf_ram.memory\[84\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10698__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07886__A2 _03652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05441__S0 _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10841_ _01210_ io_in[4] u_cpu.rf_ram.memory\[104\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09990__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10772_ _01141_ io_in[4] u_cpu.rf_ram.memory\[95\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07638__A2 _03513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05649__A1 _01490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06310__A2 _02745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__04872__A2 _01443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09260__A1 _04448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08063__A2 _03760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10078__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07810__A2 u_cpu.cpu.state.o_cnt_r\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05821__A1 _01467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09012__A1 _04434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10206_ _00592_ io_in[4] u_cpu.rf_ram.memory\[14\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09563__A2 _04762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06377__A2 _02784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10137_ _00523_ io_in[4] u_cpu.rf_ram.memory\[142\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05517__B _01534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09315__A2 _04613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10068_ _00462_ io_in[4] u_cpu.rf_ram.memory\[56\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07877__A2 _03652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05432__S0 _01530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06301__A2 _02733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06230_ _02669_ _02697_ _02698_ _00112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04863__A2 u_cpu.cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09713__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06161_ _02628_ _02642_ _02643_ _00098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08054__A2 _03750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05112_ u_cpu.rf_ram.memory\[124\]\[1\] u_cpu.rf_ram.memory\[125\]\[1\] u_cpu.rf_ram.memory\[126\]\[1\]
+ u_cpu.rf_ram.memory\[127\]\[1\] _01496_ _01594_ _01696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_06092_ _02402_ u_scanchain_local.module_data_in\[68\] _02478_ u_arbiter.i_wb_cpu_dbus_adr\[31\]
+ _02583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07801__A2 _03605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09920_ _00314_ io_in[4] u_cpu.rf_ram.memory\[77\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05812__A1 _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05043_ _01621_ _01627_ _01628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09863__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09554__A2 _04762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09851_ _00245_ io_in[4] u_cpu.rf_ram.memory\[50\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06368__A2 u_cpu.cpu.immdec.imm11_7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07565__A1 _03318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08802_ u_cpu.cpu.ctrl.o_ibus_adr\[9\] _04309_ _04311_ u_cpu.cpu.ctrl.o_ibus_adr\[10\]
+ _04321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_112_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09782_ _00176_ io_in[4] u_cpu.rf_ram.memory\[46\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06994_ u_cpu.rf_ram.memory\[60\]\[3\] _03147_ _03151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10840__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08733_ _04279_ _01035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09306__A2 _04613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05945_ _02464_ _02465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07317__A1 _03322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08664_ _03703_ _04237_ _04243_ _01002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05876_ u_arbiter.i_wb_cpu_rdt\[9\] u_arbiter.i_wb_cpu_dbus_dat\[6\] _02418_ _02424_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07615_ u_cpu.rf_ram.memory\[22\]\[2\] _03496_ _03501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05423__S0 _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08595_ _03909_ _04185_ _04186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10990__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07546_ u_cpu.rf_ram.memory\[132\]\[5\] _03455_ _03461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08293__A2 u_arbiter.i_wb_cpu_rdt\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07477_ _03320_ _03415_ _03422_ _00635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10220__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09216_ _04440_ _04563_ _04566_ _01231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06428_ u_cpu.rf_ram.memory\[44\]\[0\] _02816_ _02817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09147_ u_cpu.rf_ram.memory\[103\]\[4\] _04523_ _04528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09242__A1 _04448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06359_ _02687_ _02770_ _02775_ _00164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08045__A2 _03750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09078_ _04490_ _01169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10370__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05803__A1 _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08029_ u_cpu.rf_ram.memory\[11\]\[2\] _03740_ _03743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11040_ _01409_ io_in[4] u_cpu.rf_ram.memory\[100\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09545__A2 _04752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06359__A2 _02770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05031__A2 _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08505__B1 _04106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06531__A2 _02872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10824_ _01193_ io_in[4] u_cpu.rf_ram.memory\[102\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05072__B _01519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10755_ _01124_ io_in[4] u_cpu.rf_ram.memory\[97\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09736__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10686_ _01056_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10713__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08036__A2 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09886__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07795__A1 _02395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10863__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09536__A2 _04752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07547__A1 _03318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08347__I0 u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06770__A2 _03018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05730_ _01445_ _02305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05661_ u_cpu.rf_ram.memory\[68\]\[7\] u_cpu.rf_ram.memory\[69\]\[7\] u_cpu.rf_ram.memory\[70\]\[7\]
+ u_cpu.rf_ram.memory\[71\]\[7\] _01507_ _01605_ _02239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_90_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06522__A2 _02870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10243__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07400_ u_cpu.rf_ram.memory\[138\]\[4\] _03375_ _03380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08380_ _03999_ _04001_ _03969_ _04002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_1_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05592_ _01473_ _02121_ _02170_ _00006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_17_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07331_ _03318_ _03335_ _03341_ _00570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09472__A1 _04622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08275__A2 _02411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06286__A1 u_cpu.cpu.immdec.imm11_7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07262_ u_cpu.rf_ram.memory\[13\]\[2\] _03297_ _03300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09001_ u_cpu.rf_ram.memory\[94\]\[5\] _04436_ _04447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10393__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06213_ _02685_ _02679_ _02686_ _00107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05884__I1 u_arbiter.i_wb_cpu_dbus_dat\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09224__A1 _04448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08027__A2 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07193_ _02647_ _03257_ _03261_ _00512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06144_ u_cpu.rf_ram_if.wdata1_r\[0\] _02606_ _02629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__06589__A2 _02285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06075_ _02403_ _02566_ _02568_ _02569_ _00087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_28_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05026_ u_cpu.rf_ram.memory\[92\]\[0\] u_cpu.rf_ram.memory\[93\]\[0\] u_cpu.rf_ram.memory\[94\]\[0\]
+ u_cpu.rf_ram.memory\[95\]\[0\] _01562_ _01563_ _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09903_ _00297_ io_in[4] u_cpu.rf_ram.memory\[129\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09834_ _00228_ io_in[4] u_cpu.rf_ram.memory\[48\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06210__A1 _02683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05872__S _02418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05644__S0 _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08750__A3 _02598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09765_ _00159_ io_in[4] u_cpu.rf_ram.memory\[80\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06977_ _03106_ _03137_ _03141_ _00416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_73_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06761__A2 _02814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08468__B _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08716_ u_arbiter.i_wb_cpu_dbus_adr\[15\] u_arbiter.i_wb_cpu_dbus_adr\[16\] _04257_
+ _04271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_73_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05928_ _02450_ _02403_ _02451_ _00055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09696_ _04844_ _01433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_73_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08647_ u_cpu.cpu.genblk3.csr.timer_irq_r _04233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_54_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05859_ u_arbiter.i_wb_cpu_rdt\[2\] _02414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09759__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05316__A3 _01897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06513__A2 _02861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08578_ u_cpu.cpu.immdec.imm19_12_20\[3\] _04171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_70_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07529_ _03318_ _03445_ _03451_ _00658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10736__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08266__A2 u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10540_ _00913_ io_in[4] u_cpu.rf_ram.memory\[33\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10471_ _00844_ io_in[4] u_cpu.rf_ram.memory\[118\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08018__A2 _03730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06029__A1 _02461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10886__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10116__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07529__A1 _03318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11023_ _01392_ io_in[4] u_cpu.rf_ram.memory\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06201__A1 _02675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05635__S0 _01529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06752__A2 _03008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10266__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07701__A1 _03508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10807_ _01176_ io_in[4] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09454__A1 _04622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08257__A2 _03885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06268__A1 _02669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05530__B _01558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10738_ _01107_ io_in[4] u_cpu.rf_ram.memory\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09206__A1 _04448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05866__I1 u_arbiter.i_wb_cpu_dbus_dat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08009__A2 _03730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10669_ _01042_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08414__C1 _03988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08560__C _04031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05779__B1 _02291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05756__I _02330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11041__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06900_ u_cpu.rf_ram.memory\[64\]\[5\] _03089_ _03095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06991__A2 _03147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07880_ _03502_ _03652_ _03656_ _00805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10609__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08193__A1 u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05626__S0 _01576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06831_ _02895_ _03049_ _03056_ _00355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06743__A2 _02780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07940__A1 _03508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09901__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09550_ u_cpu.rf_ram.memory\[26\]\[1\] _04762_ _04764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06762_ _03017_ _03018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_48_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08501_ _03955_ _04101_ _04104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05713_ _01447_ _01449_ _02289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10759__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09481_ u_cpu.rf_ram.memory\[88\]\[5\] _04711_ _04717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09693__A1 _02273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06693_ u_cpu.rf_ram.memory\[129\]\[1\] _02978_ _02980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08432_ _03699_ _04041_ _04045_ _00968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05644_ u_cpu.rf_ram.memory\[112\]\[7\] u_cpu.rf_ram.memory\[113\]\[7\] u_cpu.rf_ram.memory\[114\]\[7\]
+ u_cpu.rf_ram.memory\[115\]\[7\] _01572_ _01573_ _02222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_91_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08363_ _03914_ _03903_ _03986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08248__A2 _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05575_ u_cpu.rf_ram.memory\[72\]\[6\] u_cpu.rf_ram.memory\[73\]\[6\] u_cpu.rf_ram.memory\[74\]\[6\]
+ u_cpu.rf_ram.memory\[75\]\[6\] _01562_ _01563_ _02154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07314_ u_cpu.rf_ram.memory\[73\]\[6\] _03325_ _03332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08294_ _02464_ _03920_ _03921_ _03922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07245_ _03104_ _03287_ _03290_ _00535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05482__A2 _02057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07176_ u_cpu.rf_ram.memory\[9\]\[4\] _03247_ _03252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10139__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08956__B1 _03969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06127_ u_cpu.cpu.immdec.imm11_7\[1\] _02611_ _02612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06431__A1 _02681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06058_ _02555_ _02548_ _02397_ _02556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_78_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06982__A2 _03137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10289__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05009_ _01499_ _01594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08184__A1 u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05617__S0 _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08184__B2 u_arbiter.i_wb_cpu_dbus_dat\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09817_ _00211_ io_in[4] u_cpu.rf_ram.memory\[41\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06734__A2 _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09748_ _00142_ io_in[4] u_cpu.rf_ram.memory\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09679_ _04628_ _04832_ _04835_ _01425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06498__A1 _02689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08645__C _04231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09436__A1 _04622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08239__A2 _03808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05170__A1 _01746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05350__B _01518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07998__A1 _03701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10523_ _00896_ io_in[4] u_cpu.rf_ram.memory\[115\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06670__A1 _02743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05473__A2 _02043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10454_ _00827_ io_in[4] u_cpu.rf_ram.memory\[117\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11064__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08947__B1 _03962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08411__A2 _03956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10385_ _00758_ io_in[4] u_cpu.rf_ram.memory\[37\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06422__A1 _02691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06973__A2 _03137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09924__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08175__A1 u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11006_ _01375_ io_in[4] u_cpu.rf_ram.memory\[25\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05608__S0 _01530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06725__A2 _02803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07922__A1 _03508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10901__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06200__I _02676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09675__A1 _04622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08478__A2 _04075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07150__A2 _03237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05360_ u_cpu.rf_ram.memory\[52\]\[4\] u_cpu.rf_ram.memory\[53\]\[4\] u_cpu.rf_ram.memory\[54\]\[4\]
+ u_cpu.rf_ram.memory\[55\]\[4\] _01572_ _01573_ _01941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_14_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05291_ _01597_ _01872_ _01600_ _01873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07966__I _02666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07030_ u_cpu.rf_ram.memory\[5\]\[3\] _03167_ _03171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08402__A2 _03988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10431__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08981_ u_cpu.rf_ram.memory\[97\]\[7\] _04425_ _04433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06964__A2 _03127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07932_ _03500_ _03682_ _03685_ _00828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08166__A1 u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07863_ _03642_ _03643_ _03645_ _02348_ _03646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10581__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06716__A2 _02988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06814_ u_cpu.rf_ram.memory\[6\]\[7\] _03039_ _03047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09602_ u_cpu.rf_ram.memory\[0\]\[0\] _04792_ _04793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07794_ _02263_ _02914_ _03602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09533_ _04626_ _04752_ _04754_ _01360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06745_ u_cpu.rf_ram.memory\[74\]\[0\] _03008_ _03009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08469__A2 _04069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09464_ _04634_ _04701_ _04707_ _01338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06676_ u_cpu.rf_ram.memory\[119\]\[2\] _02967_ _02970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07141__A2 _03227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08415_ _03935_ _03976_ _04033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_12_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05627_ _01597_ _02204_ _01579_ _02205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09395_ u_cpu.rf_ram.memory\[85\]\[7\] _04661_ _04669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09418__A1 _04622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05152__A1 _01473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08346_ _03922_ _03923_ _03971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05558_ u_cpu.rf_ram.memory\[116\]\[6\] u_cpu.rf_ram.memory\[117\]\[6\] u_cpu.rf_ram.memory\[118\]\[6\]
+ u_cpu.rf_ram.memory\[119\]\[6\] _01576_ _01577_ _02137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_138_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08277_ u_arbiter.i_wb_cpu_rdt\[14\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[14\]
+ _02465_ _03905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05489_ u_cpu.rf_ram.memory\[76\]\[5\] u_cpu.rf_ram.memory\[77\]\[5\] u_cpu.rf_ram.memory\[78\]\[5\]
+ u_cpu.rf_ram.memory\[79\]\[5\] _01529_ _01500_ _02069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08641__A2 _04165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09069__S _04485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07228_ u_cpu.rf_ram.memory\[141\]\[3\] _03277_ _03281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09947__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07159_ _03108_ _03237_ _03242_ _00497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10170_ _00556_ io_in[4] u_cpu.rf_ram.memory\[72\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10924__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06955__A2 _03127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06707__A2 _02976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07904__A1 _03508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05345__B _01482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07380__A2 _03365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05391__A1 _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09657__A1 _04622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05781__I3 u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09331__I _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07132__A2 _03227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10304__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05143__A1 _01465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08880__A2 _04361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06891__A1 _02881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08632__A2 _04218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10454__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10506_ _00879_ io_in[4] u_cpu.rf_ram.memory\[112\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06643__A1 _02891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10437_ _00810_ io_in[4] u_cpu.rf_ram.memory\[35\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08396__A1 _03910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07199__A2 _03257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10368_ _00741_ io_in[4] u_cpu.rf_ram.memory\[123\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06946__A2 _03117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10299_ _00685_ io_in[4] u_cpu.rf_ram.memory\[12\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_04860_ _01443_ _01446_ _01447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07371__A2 _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06530_ u_cpu.rf_ram.memory\[47\]\[3\] _02872_ _02876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07123__A2 _03217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05134__A1 _01617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06461_ u_cpu.rf_ram.memory\[51\]\[6\] _02829_ _02836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08871__A2 _04351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08200_ _03852_ _03853_ _00928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05412_ u_cpu.rf_ram.memory\[132\]\[4\] u_cpu.rf_ram.memory\[133\]\[4\] u_cpu.rf_ram.memory\[134\]\[4\]
+ u_cpu.rf_ram.memory\[135\]\[4\] _01641_ _01642_ _01993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09180_ _04440_ _04543_ _04546_ _01215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06392_ u_cpu.rf_ram.memory\[46\]\[1\] _02794_ _02796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08131_ u_cpu.cpu.mem_bytecnt\[1\] _02355_ _02306_ _02291_ _03799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_18_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05343_ _01528_ _01923_ _01924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08062_ _03691_ _03760_ _03761_ _00882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05274_ u_cpu.rf_ram.memory\[48\]\[3\] u_cpu.rf_ram.memory\[49\]\[3\] u_cpu.rf_ram.memory\[50\]\[3\]
+ u_cpu.rf_ram.memory\[51\]\[3\] _01576_ _01577_ _01856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10947__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07013_ _03106_ _03157_ _03161_ _00432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05988__A3 _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08387__A1 _03956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06937__A2 _03117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08964_ _02621_ _04391_ _04422_ _04423_ _01122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_102_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09416__I _04680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07915_ u_cpu.rf_ram.memory\[34\]\[3\] _03672_ _03676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08895_ _02637_ _04371_ _04373_ _01103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_97_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07846_ _03506_ _03626_ _03632_ _00794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05165__B _01534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05880__S _02418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07362__A2 _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10327__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09639__A1 _04622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07777_ _03592_ _03593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04989_ u_cpu.rf_ram.memory\[52\]\[0\] u_cpu.rf_ram.memory\[53\]\[0\] u_cpu.rf_ram.memory\[54\]\[0\]
+ u_cpu.rf_ram.memory\[55\]\[0\] _01572_ _01573_ _01574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_71_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06728_ _02881_ _02998_ _02999_ _00309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09516_ _02293_ _03605_ _04742_ _04743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_25_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08311__A1 _03901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07114__A2 _03217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09447_ u_cpu.rf_ram.memory\[111\]\[6\] _04691_ _04698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05125__A1 _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06659_ u_cpu.rf_ram.memory\[40\]\[3\] _02956_ _02960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08862__A2 _04351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10477__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06873__A1 _02881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09378_ _02667_ _04651_ _04659_ _01300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05920__I0 u_arbiter.i_wb_cpu_rdt\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08329_ _02911_ _03955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06625__A1 _02891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10222_ _00608_ io_in[4] u_cpu.rf_ram.memory\[39\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06928__A2 _03100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10153_ _00539_ io_in[4] u_cpu.rf_ram.memory\[140\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11102__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10084_ _00478_ io_in[4] u_cpu.rf_ram.memory\[54\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08550__A1 _04141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07353__A2 _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05364__B2 _01944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10986_ _01355_ io_in[4] u_cpu.cpu.genblk3.csr.mie_mtie vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08302__A1 _03917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07105__A2 _03207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05522__C _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05911__I0 u_arbiter.i_wb_cpu_rdt\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08369__A1 _03935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08369__B2 _03986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09030__A2 _04463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06919__A2 _03100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07592__A2 _03485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05961_ _02401_ _02461_ _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07700_ u_cpu.rf_ram.memory\[125\]\[6\] _03543_ _03550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04912_ _01496_ _01497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08680_ _03701_ _04247_ _04252_ _01009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05892_ _02432_ _00036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_93_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07344__A2 _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08541__A1 _03932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07631_ _03510_ _03496_ _03511_ _00700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07562_ u_cpu.rf_ram.memory\[131\]\[4\] _03465_ _03470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05450__S1 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09301_ u_cpu.rf_ram.memory\[69\]\[0\] _04613_ _04614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06513_ u_cpu.rf_ram.memory\[48\]\[4\] _02861_ _02866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09792__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07493_ _03318_ _03425_ _03431_ _00642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08844__A2 _04327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09232_ _04438_ _04573_ _04575_ _01238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05202__S1 _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06855__A1 _02881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06444_ _02614_ _02742_ _02825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_107_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09163_ u_cpu.rf_ram.memory\[104\]\[3\] _04533_ _04537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06375_ _02681_ _02784_ _02786_ _00169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__04961__S0 _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08114_ _03789_ _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05326_ _01901_ _01903_ _01905_ _01907_ _01466_ _01908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_119_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09094_ _04498_ _01177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08045_ u_cpu.rf_ram.memory\[112\]\[1\] _03750_ _03752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05257_ _01513_ _01838_ _01482_ _01839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11125__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05830__A2 _02389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09021__A2 _04453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05188_ _01764_ _01766_ _01768_ _01770_ _01581_ _01771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_118_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04999__B _01583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09996_ _00390_ io_in[4] u_cpu.rf_ram.memory\[29\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08780__A1 _02259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07583__A2 _03475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08947_ _03958_ _03947_ _04031_ _03962_ _04408_ _04409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__05594__A1 _01513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08878_ u_cpu.rf_ram.memory\[3\]\[2\] _04361_ _04364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07335__A2 _03335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07829_ u_cpu.rf_ram.memory\[91\]\[6\] _03616_ _03623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10840_ _01209_ io_in[4] u_cpu.rf_ram.memory\[104\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05623__B _01480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05441__S1 _01531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07099__A1 _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10771_ _01140_ io_in[4] u_cpu.rf_ram.memory\[95\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05649__A2 _02217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08599__A1 _03932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09260__A2 _04583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06074__A2 _02397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07271__A1 _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05821__A2 _02373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09012__A2 _04453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10205_ _00591_ io_in[4] u_cpu.rf_ram.memory\[14\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08220__B1 _03829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08771__A1 _03699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07574__A2 _03475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10136_ _00522_ io_in[4] u_cpu.rf_ram.memory\[142\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05585__A1 _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10067_ _00461_ io_in[4] u_cpu.rf_ram.memory\[56\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10642__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08523__A1 _03966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07326__A2 _03335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04928__I _01512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05432__S1 _01532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10792__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10969_ _01338_ io_in[4] u_cpu.rf_ram.memory\[87\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08826__A2 _04327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06837__A1 _02881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10022__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11148__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06160_ u_cpu.rf_ram.memory\[82\]\[2\] _02628_ _02643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__04863__A3 _01442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09251__A2 _04583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05111_ _01688_ _01690_ _01692_ _01694_ _01560_ _01695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_06091_ u_cpu.cpu.ctrl.o_ibus_adr\[31\] _02578_ _02582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_102_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05042_ u_cpu.rf_ram.memory\[72\]\[0\] u_cpu.rf_ram.memory\[73\]\[0\] u_cpu.rf_ram.memory\[74\]\[0\]
+ u_cpu.rf_ram.memory\[75\]\[0\] _01522_ _01622_ _01627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_144_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10172__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08211__B1 _03833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09850_ _00244_ io_in[4] u_cpu.rf_ram.memory\[50\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08762__A1 _02677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06368__A3 _02622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07565__A2 _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08801_ _04320_ _01062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_140_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05576__A1 _01621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06993_ _03104_ _03147_ _03150_ _00423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09781_ _00175_ io_in[4] u_cpu.rf_ram.memory\[42\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05944_ u_cpu.cpu.genblk1.align.ctrl_misal _02464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08732_ u_arbiter.i_wb_cpu_dbus_adr\[23\] u_arbiter.i_wb_cpu_dbus_adr\[24\] _02335_
+ _04279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08514__A1 _04111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07317__A2 _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08514__B2 _03910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05328__A1 _01473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08663_ u_cpu.rf_ram.memory\[32\]\[5\] _04237_ _04243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05875_ _02423_ _00028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_81_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05423__S1 _01509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07614_ _02641_ _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08594_ u_arbiter.i_wb_cpu_rdt\[16\] u_arbiter.i_wb_cpu_rdt\[0\] _02466_ _04185_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07545_ _03316_ _03455_ _03460_ _00665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08754__B _02292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07476_ u_cpu.rf_ram.memory\[136\]\[6\] _03415_ _03422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09215_ u_cpu.rf_ram.memory\[105\]\[2\] _04563_ _04566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06427_ _02815_ _02816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09146_ _04442_ _04523_ _04527_ _01200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06358_ u_cpu.rf_ram.memory\[78\]\[4\] _02770_ _02775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09242__A2 _04573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10515__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05309_ u_cpu.rf_ram.memory\[68\]\[3\] u_cpu.rf_ram.memory\[69\]\[3\] u_cpu.rf_ram.memory\[70\]\[3\]
+ u_cpu.rf_ram.memory\[71\]\[3\] _01507_ _01605_ _01891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07253__A1 _03112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09077_ u_arbiter.i_wb_cpu_rdt\[20\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[4\]
+ _04485_ _04490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06289_ u_cpu.rf_ram.memory\[1\]\[0\] _02733_ _02734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09077__S _04485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08028_ _02637_ _03740_ _03742_ _00867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05654__I2 u_cpu.rf_ram.memory\[82\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08202__B1 _03833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05618__B _01558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10665__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07556__A2 _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05567__A1 _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05337__C _01486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09979_ _00373_ io_in[4] u_cpu.rf_ram.memory\[65\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07308__A2 _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05319__A1 _01465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10823_ _01192_ io_in[4] u_cpu.rf_ram.memory\[102\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08808__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10045__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06819__A1 _02881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10754_ _01123_ io_in[4] u_cpu.rf_ram.memory\[97\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09481__A2 _04711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06295__A2 _02733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10685_ _01055_ io_in[4] u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04925__S0 _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09233__A2 _04573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10195__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07547__A2 _03455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10119_ _00513_ io_in[4] u_cpu.rf_ram.memory\[15\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11099_ _00028_ io_in[0] u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05660_ _01621_ _02237_ _02238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05591_ _02160_ _02169_ _02170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07330_ u_cpu.rf_ram.memory\[71\]\[5\] _03335_ _03341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09472__A2 _04711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10538__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07483__A1 _03306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07261_ _02637_ _03297_ _03299_ _00542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06286__A2 _02622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09000_ _02656_ _04446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06212_ u_cpu.rf_ram.memory\[21\]\[3\] _02679_ _02686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07192_ u_cpu.rf_ram.memory\[15\]\[3\] _03257_ _03261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09830__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09224__A2 _04563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07235__A1 _03112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06143_ _02627_ _02628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10688__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07786__A2 _03593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06074_ u_arbiter.i_wb_cpu_dbus_adr\[27\] _02397_ _02402_ _02569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_133_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05797__A1 _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05025_ _01490_ _01593_ _01609_ _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_09902_ _00296_ io_in[4] u_cpu.rf_ram.memory\[129\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09980__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05438__B _01518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07538__A2 _03455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09833_ _00227_ io_in[4] u_cpu.rf_ram.memory\[48\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06210__A2 _02679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05644__S1 _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09764_ _00158_ io_in[4] u_cpu.rf_ram.memory\[80\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06976_ u_cpu.rf_ram.memory\[61\]\[3\] _03137_ _03141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08715_ _04270_ _01026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05927_ _02403_ u_scanchain_local.module_data_in\[35\] _02451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09695_ _02273_ u_cpu.rf_ram.rdata\[7\] u_cpu.rf_ram_if.rtrig0 _04844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_66_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10068__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09160__A1 _04438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08646_ _04232_ _00995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_05858_ _02411_ _02403_ _02413_ _02408_ _00070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_70_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07710__A2 _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_55_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08577_ _04169_ _04165_ _04170_ _04003_ _00988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05789_ _02361_ _02362_ _02363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07528_ u_cpu.rf_ram.memory\[133\]\[5\] _03445_ _03451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09463__A2 _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06277__A2 _02719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07459_ _03320_ _03405_ _03412_ _00627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10470_ _00843_ io_in[4] u_cpu.rf_ram.memory\[118\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08704__S _04257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09215__A2 _04563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09129_ u_cpu.rf_ram.memory\[102\]\[4\] _04513_ _04518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08974__A1 _03699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07529__A2 _03445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11022_ _01391_ io_in[4] u_cpu.rf_ram.memory\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06201__A2 _02677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05635__S1 _01500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09334__I _02656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09703__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05399__S0 _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07701__A2 _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05712__A1 _01441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10806_ _01175_ io_in[4] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09454__A2 _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09853__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06268__A2 _02719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07465__A1 _03306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10737_ _01106_ io_in[4] u_cpu.rf_ram.memory\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10830__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09206__A2 _04553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05571__S0 _01522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10668_ _01041_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07217__A1 _03112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08414__B1 _03909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10599_ _00972_ io_in[4] u_cpu.rf_ram.memory\[114\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08414__C2 _03945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08965__A1 _02695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07768__A2 _03583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05779__A1 _02285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10980__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06440__A2 _02816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09390__A1 _04632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08193__A2 _03822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05626__S1 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06830_ u_cpu.rf_ram.memory\[68\]\[6\] _03049_ _03056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10210__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07940__A2 _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06761_ _02768_ _02814_ _03017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05951__A1 _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09142__A1 _04438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08500_ u_cpu.cpu.immdec.imm30_25\[1\] _03956_ _03959_ _04099_ _04102_ _04103_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_23_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05712_ _01441_ _02284_ _02286_ _02288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09480_ _04632_ _04711_ _04716_ _01345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06692_ _02881_ _02978_ _02979_ _00293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09693__A2 _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08431_ u_cpu.rf_ram.memory\[114\]\[3\] _04041_ _04045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05643_ _01566_ _02220_ _01558_ _02221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10360__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08362_ _03974_ _03908_ _03985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05574_ _01617_ _02152_ _01519_ _02153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09445__A2 _04691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07313_ _03318_ _03325_ _03331_ _00562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07456__A1 u_cpu.rf_ram.memory\[49\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06259__A2 _02707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08293_ _02464_ u_arbiter.i_wb_cpu_rdt\[11\] _03921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07244_ u_cpu.rf_ram.memory\[140\]\[2\] _03287_ _03290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05562__S0 _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05012__I _01504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07175_ _02647_ _03247_ _03251_ _00504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05947__I _02466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08956__A1 _03947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06126_ _02606_ _02611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__04851__I _01438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06431__A2 _02816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06057_ u_cpu.cpu.ctrl.o_ibus_adr\[24\] _02555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_114_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05008_ _01586_ _01588_ _01590_ _01592_ _01560_ _01593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_8_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09726__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08184__A2 _03822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09816_ _00210_ io_in[4] u_cpu.rf_ram.memory\[41\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05617__S1 _01531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07931__A2 _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09747_ _00141_ io_in[4] u_cpu.rf_ram.memory\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05942__A1 _02388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10703__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06959_ _03106_ _03127_ _03131_ _00408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09678_ u_cpu.rf_ram.memory\[23\]\[2\] _04832_ _04835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09684__A2 _04832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09876__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07695__A1 _03502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08629_ _03896_ _04215_ _04217_ _04218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06498__A2 _02851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10853__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09436__A2 _04691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05170__A2 _01748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07447__A1 _03306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07998__A2 _03720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10522_ _00895_ io_in[4] u_cpu.rf_ram.memory\[115\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10453_ _00826_ io_in[4] u_cpu.rf_ram.memory\[117\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05473__A3 _02052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06670__A2 _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08947__A1 _03958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10384_ _00757_ io_in[4] u_cpu.rf_ram.memory\[37\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06422__A2 _02805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10233__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09372__A1 _02652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08175__A2 _03822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11005_ _01374_ io_in[4] u_cpu.rf_ram.memory\[26\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05608__S1 _01532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07922__A2 _03672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10383__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09124__A1 _04438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09675__A2 _04832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07686__A1 _02803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06489__A2 _02851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09427__A2 _04681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07989__A2 _03720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05290_ u_cpu.rf_ram.memory\[120\]\[3\] u_cpu.rf_ram.memory\[121\]\[3\] u_cpu.rf_ram.memory\[122\]\[3\]
+ u_cpu.rf_ram.memory\[123\]\[3\] _01598_ _01556_ _01872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06110__A1 _02259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06661__A2 _02956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08938__A1 _02728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09749__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07610__A1 _03494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06413__A2 _02805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08980_ _03705_ _04425_ _04432_ _01129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07931_ u_cpu.rf_ram.memory\[117\]\[2\] _03682_ _03685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10726__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08166__A2 _02915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07862_ _03644_ _02334_ _01441_ _01442_ _03645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_112_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09899__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09601_ _04791_ _04792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07913__A2 _03672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06813_ _02662_ _03039_ _03046_ _00347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_110_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07793_ _03510_ _03593_ _03601_ _00772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09532_ u_cpu.rf_ram.memory\[27\]\[1\] _04752_ _04754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06744_ _03007_ _03008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10876__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09666__A2 _04822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09463_ u_cpu.rf_ram.memory\[87\]\[5\] _04701_ _04707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07677__A1 _03502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06675_ _02885_ _02967_ _02969_ _00286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08414_ _03940_ _03908_ _03909_ _04030_ _03988_ _03945_ _04032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__05451__B _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05626_ u_cpu.rf_ram.memory\[48\]\[7\] u_cpu.rf_ram.memory\[49\]\[7\] u_cpu.rf_ram.memory\[50\]\[7\]
+ u_cpu.rf_ram.memory\[51\]\[7\] _01576_ _01577_ _02204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09394_ _04636_ _04661_ _04668_ _01307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09418__A2 _04681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10106__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07429__A1 _03306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05557_ _01602_ _02135_ _02136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08345_ _03909_ _03917_ _03970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05170__C _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05878__S _02418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08276_ _03901_ _03903_ _03904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06101__A1 u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05488_ _01621_ _02067_ _02068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07227_ _03104_ _03277_ _03280_ _00527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10256__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08929__A1 _02264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08929__B2 _04160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07158_ u_cpu.rf_ram.memory\[52\]\[4\] _03237_ _03242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06109_ _02307_ _02311_ _02598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06404__A2 _02794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07601__A1 _02657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08988__I _02636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07089_ _03110_ _03197_ _03203_ _00466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09085__S _04485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09354__A1 _04632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08401__I0 u_arbiter.i_wb_cpu_rdt\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06168__A1 _02606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07904__A2 _03662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09106__A1 _04438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05230__I3 u_cpu.rf_ram.memory\[139\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09657__A2 _04822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05391__A2 _01971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07668__A1 _02766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09409__A2 _04671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11031__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06891__A2 _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08617__B1 _03909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08391__C _03938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10505_ _00878_ io_in[4] u_cpu.rf_ram.memory\[112\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07840__A1 _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06643__A2 _02945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10436_ _00809_ io_in[4] u_cpu.rf_ram.memory\[92\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10749__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09593__A1 _04632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10367_ _00014_ io_in[4] u_cpu.rf_ram_if.rdata0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10298_ _00684_ io_in[4] u_cpu.rf_ram.memory\[130\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__04957__A2 _01535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08148__A2 _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10899__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06211__I _02646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09648__A2 _04812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10129__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07659__A1 _03502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08320__A2 _03947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05271__B _01480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06460_ _02689_ _02829_ _02835_ _00205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06331__A1 _02681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05411_ _01465_ _01991_ _01992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06391_ _02669_ _02794_ _02795_ _00176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06882__A2 _03079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10279__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08130_ _03707_ _03790_ _03798_ _00913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05342_ u_cpu.rf_ram.memory\[8\]\[4\] u_cpu.rf_ram.memory\[9\]\[4\] u_cpu.rf_ram.memory\[10\]\[4\]
+ u_cpu.rf_ram.memory\[11\]\[4\] _01523_ _01525_ _01923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08084__A1 _03697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08061_ u_cpu.rf_ram.memory\[122\]\[0\] _03760_ _03761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06634__A2 _02945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05273_ _01571_ _01854_ _01855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07012_ u_cpu.rf_ram.memory\[19\]\[3\] _03157_ _03161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08963_ u_cpu.cpu.immdec.imm30_25\[0\] _03897_ _04391_ _04423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_142_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05070__A1 _01513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09336__A1 _04634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07914_ _03500_ _03672_ _03675_ _00820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08894_ u_cpu.rf_ram.memory\[2\]\[1\] _04371_ _04373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07845_ u_cpu.rf_ram.memory\[90\]\[5\] _03626_ _03632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07898__A1 _03502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07776_ _02717_ _02782_ _03592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09639__A2 _04812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04988_ _01499_ _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08476__C _04031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09515_ u_cpu.cpu.decode.co_ebreak u_cpu.cpu.mem_bytecnt\[1\] _02291_ _02290_ _04742_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__11054__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06727_ u_cpu.rf_ram.memory\[77\]\[0\] _02998_ _02999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08311__A2 _03938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09446_ _04634_ _04691_ _04697_ _01330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06322__A1 _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06658_ _02887_ _02956_ _02959_ _00279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05609_ _01464_ _02186_ _01481_ _02187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06873__A2 _03079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09377_ u_cpu.rf_ram.memory\[10\]\[7\] _04651_ _04659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06589_ _01444_ _02285_ _02913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09914__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08328_ _02328_ _03897_ _03954_ _00955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_20_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07822__A1 _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06625__A2 _02935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08259_ _03701_ _03885_ _03890_ _00950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08712__S _04257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09575__A1 _04632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10221_ _00607_ io_in[4] u_cpu.rf_ram.memory\[39\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10152_ _00538_ io_in[4] u_cpu.rf_ram.memory\[140\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07050__A2 _03177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09327__A1 _04628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05061__A1 _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10083_ _00477_ io_in[4] u_cpu.rf_ram.memory\[54\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07889__A1 _02782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05364__A2 _01940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08838__B1 _04329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10985_ _01354_ io_in[4] u_cpu.cpu.genblk3.csr.mstatus_mpie vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10421__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06864__A2 _03069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08066__A1 _03697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10571__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06616__A2 _02935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07813__A1 _02396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10419_ _00792_ io_in[4] u_cpu.rf_ram.memory\[90\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09318__A1 _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05052__A1 _01465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05266__B _01558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05960_ u_cpu.cpu.ctrl.o_ibus_adr\[5\] _02476_ _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11077__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04911_ _01495_ _01496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05891_ u_arbiter.i_wb_cpu_rdt\[16\] u_arbiter.i_wb_cpu_dbus_dat\[13\] _02431_ _02432_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07630_ u_cpu.rf_ram.memory\[22\]\[7\] _03496_ _03511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08541__A2 _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07561_ _03314_ _03465_ _03469_ _00672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09937__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09300_ _04612_ _04613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06512_ _02685_ _02861_ _02865_ _00227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07492_ u_cpu.rf_ram.memory\[135\]\[5\] _03425_ _03431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06304__A1 _02667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09231_ u_cpu.rf_ram.memory\[106\]\[1\] _04573_ _04575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06855__A2 _03069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06443_ _02693_ _02816_ _02824_ _00199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10914__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09162_ _04440_ _04533_ _04536_ _01207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06374_ u_cpu.rf_ram.memory\[42\]\[1\] _02784_ _02786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__04961__S1 _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05325_ _01638_ _01906_ _01534_ _01907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08113_ _02695_ _02782_ _03789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07804__A1 _02395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09093_ u_arbiter.i_wb_cpu_rdt\[28\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[12\]
+ _04485_ _04498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08044_ _03691_ _03750_ _03751_ _00874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05256_ u_cpu.rf_ram.memory\[12\]\[3\] u_cpu.rf_ram.memory\[13\]\[3\] u_cpu.rf_ram.memory\[14\]\[3\]
+ u_cpu.rf_ram.memory\[15\]\[3\] _01530_ _01532_ _01838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08532__S _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07280__A2 _03308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05020__I _01498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09557__A1 _04632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05291__A1 _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05187_ _01505_ _01769_ _01579_ _01770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_115_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07032__A2 _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09995_ _00389_ io_in[4] u_cpu.rf_ram.memory\[29\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05043__A1 _01621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08780__A2 _02598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08946_ _03940_ _03910_ _04408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05891__S _02431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08877_ _02637_ _04361_ _04363_ _01095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_57_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07828_ _03506_ _03616_ _03622_ _00786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10444__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07759_ _03582_ _03583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_44_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07099__A2 _03207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10770_ _01139_ io_in[4] u_cpu.rf_ram.memory\[95\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10594__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09429_ u_cpu.rf_ram.memory\[86\]\[6\] _04681_ _04688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05649__A3 _02226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06846__A2 _03059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08048__A1 _03697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08599__A2 _03998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07271__A2 _03297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05282__A1 _01548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05865__I _02388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09337__I _02661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10204_ _00590_ io_in[4] u_cpu.rf_ram.memory\[14\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08220__A1 u_arbiter.i_wb_cpu_rdt\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05034__A1 _01617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08771__A2 _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10135_ _00521_ io_in[4] u_cpu.rf_ram.memory\[142\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05086__B _01518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05585__A2 _02163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06782__A1 _02881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10066_ _00460_ io_in[4] u_cpu.rf_ram.memory\[57\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08523__A2 _04121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10937__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08287__A1 _03914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10968_ _01337_ io_in[4] u_cpu.rf_ram.memory\[87\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06837__A2 _03059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10899_ _01268_ io_in[4] u_cpu.rf_ram.memory\[108\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__04944__I _01494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09087__I0 u_arbiter.i_wb_cpu_rdt\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05110_ _01566_ _01693_ _01558_ _01694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_117_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06090_ _02576_ _02581_ _00090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07262__A2 _03297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10317__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05273__A1 _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09539__A1 _04632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05041_ _01617_ _01625_ _01519_ _01626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07014__A2 _03157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08211__A1 u_arbiter.i_wb_cpu_rdt\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08211__B2 u_arbiter.i_wb_cpu_dbus_dat\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05025__A1 _01490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08800_ u_cpu.cpu.ctrl.o_ibus_adr\[8\] _04309_ _04311_ u_cpu.cpu.ctrl.o_ibus_adr\[9\]
+ _04320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08762__A2 _02766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10467__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09780_ _00174_ io_in[4] u_cpu.rf_ram.memory\[42\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05576__A2 _02154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06992_ u_cpu.rf_ram.memory\[60\]\[2\] _03147_ _03150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08731_ _04278_ _01034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05943_ _02462_ _02463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08662_ _03701_ _04237_ _04242_ _01001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06525__A1 _02669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05874_ u_arbiter.i_wb_cpu_rdt\[8\] u_arbiter.i_wb_cpu_dbus_dat\[5\] _02418_ _02423_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_26_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07613_ _03498_ _03496_ _03499_ _00694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_54_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08593_ _01439_ _04165_ _04183_ _04184_ _00990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__05443__C _01560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07544_ u_cpu.rf_ram.memory\[132\]\[4\] _03455_ _03460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05015__I _01480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08754__C _02914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06828__A2 _03049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07475_ _03318_ _03415_ _03421_ _00634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09214_ _04438_ _04563_ _04565_ _01230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06426_ _02782_ _02814_ _02815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09145_ u_cpu.rf_ram.memory\[103\]\[3\] _04523_ _04527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06357_ _02685_ _02770_ _02774_ _00163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05886__S _02418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05308_ _01621_ _01889_ _01890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09076_ _04489_ _01168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07253__A2 _03287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06288_ _02732_ _02733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05264__A1 _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08027_ u_cpu.rf_ram.memory\[11\]\[1\] _03740_ _03742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05239_ _01812_ _01821_ _01822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08202__A1 u_arbiter.i_wb_cpu_rdt\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08202__B2 u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05016__A1 _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09978_ _00372_ io_in[4] u_cpu.rf_ram.memory\[66\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06764__A1 _02881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05567__A2 _02145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09093__S _04485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08929_ _02264_ _04391_ _04392_ _04160_ _01118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_131_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05634__B _01518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06516__A1 _02689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10822_ _01191_ io_in[4] u_cpu.rf_ram.memory\[102\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06819__A2 _03049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10753_ _01122_ io_in[4] u_cpu.cpu.immdec.imm11_7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05878__I0 u_arbiter.i_wb_cpu_rdt\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09069__I0 u_arbiter.i_wb_cpu_rdt\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10684_ _01054_ io_in[4] u_arbiter.i_wb_cpu_ibus_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07492__A2 _03425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04925__S1 _01509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07244__A2 _03287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05255__A1 _01528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08992__A2 _04436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05007__A1 _01566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09782__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11167_ u_scanchain_local.data_out io_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10118_ _00512_ io_in[4] u_cpu.rf_ram.memory\[15\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11098_ _00027_ io_in[0] u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04939__I _01499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10049_ _00443_ io_in[4] u_cpu.rf_ram.memory\[5\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11115__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05590_ _02162_ _02164_ _02166_ _02168_ _01466_ _02169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_51_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08347__S _02466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07260_ u_cpu.rf_ram.memory\[13\]\[1\] _03297_ _03299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08680__A1 _03701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07483__A2 _03425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05333__I2 u_cpu.rf_ram.memory\[22\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06211_ _02646_ _02685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07191_ _02642_ _03257_ _03260_ _00511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06142_ _02619_ _02626_ _02627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08432__A1 _03699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07235__A2 _03277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05246__A1 _01513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06073_ u_cpu.cpu.ctrl.o_ibus_adr\[27\] _02562_ _02567_ _02568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05024_ _01596_ _01601_ _01604_ _01608_ _01581_ _01609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_09901_ _00295_ io_in[4] u_cpu.rf_ram.memory\[129\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08196__B1 _03833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09832_ _00226_ io_in[4] u_cpu.rf_ram.memory\[48\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06746__A1 _02881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09763_ _00157_ io_in[4] u_cpu.rf_ram.memory\[80\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06975_ _03104_ _03137_ _03140_ _00415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08714_ u_arbiter.i_wb_cpu_dbus_adr\[14\] u_arbiter.i_wb_cpu_dbus_adr\[15\] _04257_
+ _04270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08499__A1 _03955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05926_ u_arbiter.i_wb_cpu_dbus_dat\[30\] _02450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05454__B _02033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09694_ _04843_ _01432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_54_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09160__A2 _04533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08645_ u_cpu.cpu.immdec.imm31 _03897_ _04009_ _04230_ _04231_ _04232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_05857_ _02412_ _02355_ _02413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07171__A1 _02637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08576_ u_cpu.cpu.immdec.imm19_12_20\[3\] _03897_ _04165_ _04170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_70_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05788_ u_cpu.cpu.ctrl.pc_plus_4_cy_r u_arbiter.i_wb_cpu_ibus_adr\[0\] _02362_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__05721__A2 u_cpu.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07527_ _03316_ _03445_ _03450_ _00657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07474__A2 _03415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07458_ u_cpu.rf_ram.memory\[49\]\[6\] _03405_ _03412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06409_ u_cpu.rf_ram.memory\[45\]\[0\] _02805_ _02806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07389_ _02667_ _03365_ _03373_ _00596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_108_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09128_ _04442_ _04513_ _04517_ _01192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10632__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08423__A1 _02619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07226__A2 _03277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05237__A1 _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08974__A2 _04425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09059_ _04442_ _04476_ _04480_ _01160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05788__A2 u_arbiter.i_wb_cpu_ibus_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06985__A1 _03114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08720__S _04257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11069__D u_cpu.rf_ram_if.wdata0_r\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10782__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08187__B1 _03833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11021_ _01390_ io_in[4] u_cpu.rf_ram.memory\[24\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05096__S0 _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11138__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10012__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09151__A2 _04523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05399__S1 _01622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10162__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10805_ _01174_ io_in[4] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10736_ _01105_ io_in[4] u_cpu.rf_ram.memory\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07465__A2 _03415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08662__A1 _03701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10667_ _01040_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05571__S1 _01622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08414__A1 _03940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07217__A2 _03267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08414__B2 _04030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10598_ _00971_ io_in[4] u_cpu.rf_ram.memory\[114\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05228__A1 _01492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08965__A2 _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05539__B _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05779__A2 u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06214__I _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05258__C _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08178__B1 _03833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06728__A1 _02881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05087__S0 _01551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09390__A2 _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05400__A1 _01621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06760_ _02897_ _03008_ _03016_ _00324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06089__C _02402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09142__A2 _04523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05711_ _02285_ _02286_ _02287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10505__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06691_ u_cpu.rf_ram.memory\[129\]\[0\] _02978_ _02979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07153__A1 _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08430_ _03697_ _04041_ _04044_ _00967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_93_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05642_ u_cpu.rf_ram.memory\[120\]\[7\] u_cpu.rf_ram.memory\[121\]\[7\] u_cpu.rf_ram.memory\[122\]\[7\]
+ u_cpu.rf_ram.memory\[123\]\[7\] _01598_ _01556_ _02220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_24_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08361_ _03915_ _03918_ _03912_ _03984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05573_ u_cpu.rf_ram.memory\[68\]\[6\] u_cpu.rf_ram.memory\[69\]\[6\] u_cpu.rf_ram.memory\[70\]\[6\]
+ u_cpu.rf_ram.memory\[71\]\[6\] _01507_ _01605_ _02152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_108_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07312_ u_cpu.rf_ram.memory\[73\]\[5\] _03325_ _03331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10655__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08292_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[11\] _03920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_32_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07456__A2 _03405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05467__A1 _01566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07243_ _03102_ _03287_ _03289_ _00534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05562__S1 _01563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08405__A1 _03947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07208__A2 _03267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07174_ u_cpu.rf_ram.memory\[9\]\[3\] _03247_ _03251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08956__A2 _04031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06125_ u_cpu.cpu.decode.op26 u_cpu.cpu.decode.co_ebreak _02606_ _02610_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_117_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06967__A1 _03114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06056_ u_cpu.cpu.ctrl.o_ibus_adr\[24\] u_cpu.cpu.ctrl.o_ibus_adr\[23\] _02546_ _02554_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_133_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05007_ _01566_ _01591_ _01558_ _01592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10035__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05078__S0 _01523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09815_ _00209_ io_in[4] u_cpu.rf_ram.memory\[41\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09381__A2 _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09746_ _00140_ io_in[4] u_cpu.rf_ram.memory\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06958_ u_cpu.rf_ram.memory\[62\]\[3\] _03127_ _03131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05942__A2 _02461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09133__A2 _04513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10185__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05909_ u_arbiter.i_wb_cpu_rdt\[25\] u_arbiter.i_wb_cpu_dbus_dat\[22\] _02431_ _02441_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09677_ _04626_ _04832_ _04834_ _01424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06889_ _03088_ _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08495__B _03966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08628_ _02467_ _02414_ _03965_ _04216_ _04217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_42_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07695__A2 _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05250__S0 _01523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08559_ _04149_ _04152_ _04155_ _03914_ _04156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07447__A2 _03405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05458__A1 _01548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05002__S0 _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10521_ _00894_ io_in[4] u_cpu.rf_ram.memory\[115\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10452_ _00825_ io_in[4] u_cpu.rf_ram.memory\[34\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08947__A2 _03947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05359__B _01480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10383_ _00756_ io_in[4] u_cpu.rf_ram.memory\[38\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05630__A1 _01492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11004_ _01373_ io_in[4] u_cpu.rf_ram.memory\[26\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05069__S0 _01497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09372__A2 _04651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10528__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07383__A1 _02652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05933__A2 _02397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09820__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09124__A2 _04513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07135__A1 _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10678__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07686__A2 _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08883__A1 _02652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05241__S0 _01497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09970__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08635__A1 _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07438__A2 _03395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05449__A1 _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10719_ _01089_ io_in[4] u_cpu.rf_ram.memory\[109\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06110__A2 _02598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10058__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06949__A1 _03114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07610__A2 _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05621__A1 _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07930_ _03498_ _03682_ _03684_ _00827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09363__A2 _04651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07861_ u_cpu.cpu.alu.cmp_r _03644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_29_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09600_ _02731_ _02754_ _04791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_110_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06812_ u_cpu.rf_ram.memory\[6\]\[6\] _03039_ _03046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07792_ u_cpu.rf_ram.memory\[36\]\[7\] _03593_ _03601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05480__S0 _01507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09531_ _04622_ _04752_ _04753_ _01359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09115__A2 _04503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06743_ _02768_ _02780_ _03007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09462_ _04632_ _04701_ _04706_ _01337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07677__A2 _03533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06674_ u_cpu.rf_ram.memory\[119\]\[1\] _02967_ _02969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08413_ _03914_ _03938_ _04031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05232__S0 _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05625_ _01571_ _02202_ _02203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09393_ u_cpu.rf_ram.memory\[85\]\[6\] _04661_ _04668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08344_ _03901_ _03938_ _03969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05556_ u_cpu.rf_ram.memory\[112\]\[6\] u_cpu.rf_ram.memory\[113\]\[6\] u_cpu.rf_ram.memory\[114\]\[6\]
+ u_cpu.rf_ram.memory\[115\]\[6\] _01572_ _01573_ _02135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08626__A1 _03974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07429__A2 _03395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08275_ _02465_ _02411_ _03902_ _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05487_ u_cpu.rf_ram.memory\[72\]\[5\] u_cpu.rf_ram.memory\[73\]\[5\] u_cpu.rf_ram.memory\[74\]\[5\]
+ u_cpu.rf_ram.memory\[75\]\[5\] _01562_ _01563_ _02067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07226_ u_cpu.rf_ram.memory\[141\]\[2\] _03277_ _03280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05860__A1 u_cpu.cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07157_ _03106_ _03237_ _03241_ _00496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06108_ u_cpu.cpu.ctrl.pc_plus_offset_cy_r _02331_ _02597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07601__A2 _03485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07088_ u_cpu.rf_ram.memory\[56\]\[5\] _03197_ _03203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05612__A1 _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06039_ u_cpu.cpu.ctrl.o_ibus_adr\[21\] _02539_ _02540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_120_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09843__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09354__A2 _04641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08401__I1 u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07365__A1 _03316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10820__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09106__A2 _04503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09729_ _00123_ io_in[4] u_cpu.rf_ram.memory\[18\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07117__A1 _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09993__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07668__A2 _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08865__A1 _03701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05679__A1 _02247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05223__S0 _01522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10970__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06340__A2 _02756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08953__B _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08617__A1 _03924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08617__B2 _04202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09290__A1 _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08093__A2 _03770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10200__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10504_ _00877_ io_in[4] u_cpu.rf_ram.memory\[112\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07840__A2 _03626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05851__A1 _01441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10435_ _00808_ io_in[4] u_cpu.rf_ram.memory\[92\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09042__A1 _04448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09593__A2 _04782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10366_ _00013_ io_in[4] u_cpu.rf_ram_if.rdata0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10350__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05603__A1 _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10297_ _00683_ io_in[4] u_cpu.rf_ram.memory\[130\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09345__A2 _04641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04947__I _01531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07659__A2 _03523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05509__I2 u_cpu.rf_ram.memory\[22\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05214__S0 _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06331__A2 _02756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05410_ u_cpu.rf_ram.memory\[128\]\[4\] u_cpu.rf_ram.memory\[129\]\[4\] u_cpu.rf_ram.memory\[130\]\[4\]
+ u_cpu.rf_ram.memory\[131\]\[4\] _01641_ _01642_ _01991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08608__A1 u_cpu.cpu.immdec.imm19_12_20\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06390_ u_cpu.rf_ram.memory\[46\]\[0\] _02794_ _02795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08582__C _04052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05341_ _01528_ _01921_ _01534_ _01922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08084__A2 _03770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09281__A1 _02814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09716__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06095__A1 _01445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08060_ _03759_ _03760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05142__I0 u_cpu.rf_ram.memory\[128\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05272_ u_cpu.rf_ram.memory\[52\]\[3\] u_cpu.rf_ram.memory\[53\]\[3\] u_cpu.rf_ram.memory\[54\]\[3\]
+ u_cpu.rf_ram.memory\[55\]\[3\] _01572_ _01573_ _01854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07831__A2 _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07011_ _03104_ _03157_ _03160_ _00431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09866__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09584__A2 _04782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06398__A2 _02794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07595__A1 _02642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08792__B1 _04311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08962_ _03956_ _03922_ _04421_ _04422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10843__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09336__A2 _04624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07913_ u_cpu.rf_ram.memory\[34\]\[2\] _03672_ _03675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08893_ _02632_ _04371_ _04372_ _01102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_68_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07347__A1 _03316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07844_ _03504_ _03626_ _03631_ _00793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07898__A2 _03662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07775_ _03510_ _03583_ _03591_ _00764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10993__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04987_ _01495_ _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06570__A2 _02900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09514_ u_cpu.cpu.genblk3.csr.mie_mtie _04741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_65_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05462__B _01558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06726_ _02997_ _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_17_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08329__I _02911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08698__I1 u_arbiter.i_wb_cpu_dbus_adr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09445_ u_cpu.rf_ram.memory\[111\]\[5\] _04691_ _04697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06657_ u_cpu.rf_ram.memory\[40\]\[2\] _02956_ _02959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06322__A2 _02745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10223__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05608_ u_cpu.rf_ram.memory\[12\]\[7\] u_cpu.rf_ram.memory\[13\]\[7\] u_cpu.rf_ram.memory\[14\]\[7\]
+ u_cpu.rf_ram.memory\[15\]\[7\] _01530_ _01532_ _02186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_33_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09376_ _02662_ _04651_ _04658_ _01299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_71_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06588_ _02395_ _02912_ _00256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08327_ _03944_ _03912_ _03915_ _03918_ _03896_ _03954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_33_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05539_ _01597_ _02117_ _01579_ _02118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08075__A2 _03760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09272__A1 _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08258_ u_cpu.rf_ram.memory\[113\]\[4\] _03885_ _03890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07822__A2 _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10373__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05833__A1 u_cpu.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07209_ _03104_ _03267_ _03270_ _00519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09024__A1 _04448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08189_ u_arbiter.i_wb_cpu_dbus_dat\[11\] _03835_ _03846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10220_ _00606_ io_in[4] u_cpu.rf_ram.memory\[39\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09575__A2 _04772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10151_ _00537_ io_in[4] u_cpu.rf_ram.memory\[140\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05061__A2 _01645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09327__A2 _04624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10082_ _00476_ io_in[4] u_cpu.rf_ram.memory\[55\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07889__A2 _02825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05444__S0 _01496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06561__A2 _02883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10984_ _01353_ io_in[4] u_cpu.cpu.genblk3.csr.mcause31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08302__A3 _03929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05091__C _01560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09739__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06313__A2 _02745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10716__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08066__A2 _03760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09263__A1 _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09889__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10866__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09566__A2 _04772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10418_ _00791_ io_in[4] u_cpu.rf_ram.memory\[90\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07577__A1 _03312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10349_ _00735_ io_in[4] u_cpu.rf_ram.memory\[124\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05052__A2 _01636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09318__A2 _02717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07329__A1 _03316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08526__C2 _03959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04910_ _01494_ _01495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_78_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05890_ _02388_ _02431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06001__A1 _02463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05435__S0 _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06552__A2 _02883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05282__B _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10246__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07560_ u_cpu.rf_ram.memory\[131\]\[3\] _03465_ _03469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06511_ u_cpu.rf_ram.memory\[48\]\[3\] _02861_ _02865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07491_ _03316_ _03425_ _03430_ _00641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07501__A1 _03306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06304__A2 _02733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09230_ _04434_ _04573_ _04574_ _01237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06442_ u_cpu.rf_ram.memory\[44\]\[7\] _02816_ _02824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10396__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09161_ u_cpu.rf_ram.memory\[104\]\[2\] _04533_ _04536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__04866__A2 _01452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09254__A1 _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08057__A2 _03750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06373_ _02669_ _02784_ _02785_ _00168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08112_ _03707_ _03780_ _03788_ _00905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05324_ u_cpu.rf_ram.memory\[140\]\[3\] u_cpu.rf_ram.memory\[141\]\[3\] u_cpu.rf_ram.memory\[142\]\[3\]
+ u_cpu.rf_ram.memory\[143\]\[3\] _01641_ _01642_ _01906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09092_ _03920_ _04485_ _04497_ _01176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06607__A3 _02929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05815__A1 _01467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08043_ u_cpu.rf_ram.memory\[112\]\[0\] _03750_ _03751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05255_ _01528_ _01836_ _01837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09557__A2 _04762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05186_ u_cpu.rf_ram.memory\[48\]\[2\] u_cpu.rf_ram.memory\[49\]\[2\] u_cpu.rf_ram.memory\[50\]\[2\]
+ u_cpu.rf_ram.memory\[51\]\[2\] _01576_ _01577_ _01769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_131_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09994_ _00388_ io_in[4] u_cpu.rf_ram.memory\[64\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09309__A2 _04613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05043__A2 _01627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06240__A1 _02689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05674__S0 _01523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11021__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08945_ _04405_ _04406_ _04179_ _04407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_131_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06791__A2 _03028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08876_ u_cpu.rf_ram.memory\[3\]\[1\] _04361_ _04363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_29_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05426__S0 _01523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07827_ u_cpu.rf_ram.memory\[91\]\[5\] _03616_ _03622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06543__A2 _02883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07740__A1 _02782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07758_ _02675_ _02782_ _03582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06709_ u_cpu.rf_ram.memory\[139\]\[0\] _02988_ _02989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10739__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07689_ _03494_ _03543_ _03544_ _00725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09493__A1 u_cpu.cpu.genblk3.csr.o_new_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09428_ _04634_ _04681_ _04687_ _01322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09359_ u_cpu.rf_ram.memory\[59\]\[7\] _04641_ _04649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08048__A2 _03750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09245__A1 _02849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10889__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08950__C _03955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05806__A1 _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09548__A2 _04762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10119__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07559__A1 _03312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10203_ _00589_ io_in[4] u_cpu.rf_ram.memory\[14\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08220__A2 _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05034__A2 _01618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05665__S0 _01529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10134_ _00520_ io_in[4] u_cpu.rf_ram.memory\[142\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06782__A2 _03028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10269__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10065_ _00459_ io_in[4] u_cpu.rf_ram.memory\[57\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05417__S0 _01497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07731__A1 _03502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06534__A2 _02872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10967_ _01336_ io_in[4] u_cpu.rf_ram.memory\[87\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09484__A1 _04636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08287__A2 _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06298__A1 _02652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10898_ _01267_ io_in[4] u_cpu.rf_ram.memory\[108\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09236__A1 _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08039__A2 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06217__I _02656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07798__A1 u_cpu.cpu.state.o_cnt_r\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09539__A2 _04752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05040_ u_cpu.rf_ram.memory\[68\]\[0\] u_cpu.rf_ram.memory\[69\]\[0\] u_cpu.rf_ram.memory\[70\]\[0\]
+ u_cpu.rf_ram.memory\[71\]\[0\] _01529_ _01500_ _01625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__05273__A2 _01854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04960__I _01499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11044__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08211__A2 _03822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06222__A1 _02691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05025__A2 _01593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05656__S0 _01507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06991_ _03102_ _03147_ _03149_ _00422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06773__A2 _03018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08730_ u_arbiter.i_wb_cpu_dbus_adr\[22\] u_arbiter.i_wb_cpu_dbus_adr\[23\] _02335_
+ _04278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09904__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05942_ _02388_ _02461_ _02462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05408__S0 _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08661_ u_cpu.rf_ram.memory\[32\]\[4\] _04237_ _04242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05873_ _02422_ _00027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07722__A1 _02849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06525__A2 _02872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07612_ u_cpu.rf_ram.memory\[22\]\[1\] _03496_ _03499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08592_ u_cpu.cpu.immdec.imm19_12_20\[5\] _03897_ _04165_ _04184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_53_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07543_ _03314_ _03455_ _03459_ _00664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07474_ u_cpu.rf_ram.memory\[136\]\[5\] _03415_ _03421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09213_ u_cpu.rf_ram.memory\[105\]\[1\] _04563_ _04565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06425_ _02716_ _02765_ _02814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09227__A1 _02780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09144_ _04440_ _04523_ _04526_ _01199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06356_ u_cpu.rf_ram.memory\[78\]\[3\] _02770_ _02774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07789__A1 _03506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05307_ u_cpu.rf_ram.memory\[64\]\[3\] u_cpu.rf_ram.memory\[65\]\[3\] u_cpu.rf_ram.memory\[66\]\[3\]
+ u_cpu.rf_ram.memory\[67\]\[3\] _01522_ _01622_ _01889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_136_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09075_ u_arbiter.i_wb_cpu_rdt\[19\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[3\]
+ _04485_ _04489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06287_ _02695_ _02731_ _02732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_68_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08450__A2 _03929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08026_ _02632_ _03740_ _03741_ _00866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05238_ _01814_ _01816_ _01818_ _01820_ _01466_ _01821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_122_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05187__B _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08202__A2 _03822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05169_ _01513_ _01751_ _01482_ _01752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_103_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10411__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06213__A1 _02685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09977_ _00371_ io_in[4] u_cpu.rf_ram.memory\[66\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06764__A2 _03018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08498__B _02392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08928_ u_cpu.cpu.immdec.imm11_7\[1\] _03897_ _04391_ _04392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_58_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08859_ _03695_ _04351_ _04353_ _01087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_18_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10561__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07713__A1 _03502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06516__A2 _02861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08718__S _04257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10821_ _01190_ io_in[4] u_cpu.rf_ram.memory\[102\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09466__A1 _04636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10752_ _01121_ io_in[4] u_cpu.cpu.immdec.imm11_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09218__A1 _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10683_ _00023_ io_in[4] u_cpu.cpu.ctrl.pc_plus_4_cy_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11067__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05255__A2 _01836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06452__A1 _02681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09927__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10091__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06204__A1 _02669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11166_ io_in[0] io_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06755__A2 _03008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10904__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10117_ _00511_ io_in[4] u_cpu.rf_ram.memory\[15\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11097_ _00095_ io_in[0] u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10048_ _00442_ io_in[4] u_cpu.rf_ram.memory\[5\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07704__A1 _02814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06507__A2 _02861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08752__I0 u_arbiter.i_wb_cpu_dbus_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07180__A2 _03247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05318__I0 u_cpu.rf_ram.memory\[128\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09209__A1 _02838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08680__A2 _04247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06210_ _02683_ _02679_ _02684_ _00106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07190_ u_cpu.rf_ram.memory\[15\]\[2\] _03257_ _03260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06141_ _02625_ _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08432__A2 _04041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10434__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05246__A2 _01827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06443__A1 _02693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06072_ u_cpu.cpu.ctrl.o_ibus_adr\[27\] _02562_ _02397_ _02567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06994__A2 _03147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05023_ _01554_ _01606_ _01607_ _01608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09900_ _00294_ io_in[4] u_cpu.rf_ram.memory\[129\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08196__A1 u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09831_ _00225_ io_in[4] u_cpu.rf_ram.memory\[48\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10584__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06746__A2 _03008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06974_ u_cpu.rf_ram.memory\[61\]\[2\] _03137_ _03140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09762_ _00156_ io_in[4] u_cpu.rf_ram.memory\[80\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08713_ _04269_ _01025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05925_ _02449_ _00054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09693_ _02273_ _02272_ u_cpu.rf_ram.rdata\[7\] _04843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__08499__A2 _04101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08644_ _04173_ _04129_ _04053_ _03896_ _04231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_82_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05856_ _02306_ _02412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_27_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08538__S _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07171__A2 _03247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08575_ u_cpu.cpu.immdec.imm19_12_20\[2\] _04169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09448__A1 _04636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05787_ u_cpu.cpu.state.o_cnt_r\[2\] u_cpu.cpu.ctrl.i_iscomp _02292_ _02360_ _02361_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07526_ u_cpu.rf_ram.memory\[133\]\[4\] _03445_ _03450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08120__A1 _03697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07457_ _03318_ _03405_ _03411_ _00626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08671__A2 _04247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05897__S _02431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06408_ _02804_ _02805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_41_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07388_ u_cpu.rf_ram.memory\[14\]\[7\] _03365_ _03373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_10_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09127_ u_cpu.rf_ram.memory\[102\]\[3\] _04513_ _04517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06339_ _02689_ _02756_ _02762_ _00157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08423__A2 _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05237__A2 _01819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09058_ u_cpu.rf_ram.memory\[28\]\[3\] _04476_ _04480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10927__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08009_ u_cpu.rf_ram.memory\[8\]\[1\] _03730_ _03732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06985__A2 _03137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08187__A1 u_arbiter.i_wb_cpu_rdt\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11020_ _01389_ io_in[4] u_cpu.rf_ram.memory\[24\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07934__A1 _03502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06737__A2 _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05096__S1 _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09687__A1 _04636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05364__C _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07162__A2 _03237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10307__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10804_ _01173_ io_in[4] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10735_ _01104_ io_in[4] u_cpu.rf_ram.memory\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08662__A2 _04237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10457__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06673__A1 _02881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10666_ _01039_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10597_ _00970_ io_in[4] u_cpu.rf_ram.memory\[114\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08414__A2 _03908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09611__A1 _02687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06976__A2 _03137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08178__A1 u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08178__B2 u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06728__A2 _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07925__A1 _02675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05555__B _01558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11149_ _00083_ io_in[0] u_scanchain_local.module_data_in\[61\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05087__S1 _01524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05710_ u_cpu.cpu.bne_or_bge _02286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_64_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06690_ _02977_ _02978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_63_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08350__A1 _03974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07153__A2 _03237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05641_ _01543_ _02218_ _02219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06900__A2 _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08360_ _03950_ _03967_ _03983_ _00958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05572_ _01621_ _02150_ _02151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08157__I _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08102__A1 _03697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07311_ _03316_ _03325_ _03330_ _00561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08291_ _03906_ _03908_ _03919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08653__A2 _04237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05467__A2 _02046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06664__A1 _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07242_ u_cpu.rf_ram.memory\[140\]\[1\] _03287_ _03289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07173_ _02642_ _03247_ _03250_ _00503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_9_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08405__A2 _03972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06416__A1 _02685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06124_ _02606_ _02607_ _02608_ _02264_ _02609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_105_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06967__A2 _03127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06055_ _02389_ u_scanchain_local.module_data_in\[61\] _02553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08169__A1 u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05006_ u_cpu.rf_ram.memory\[104\]\[0\] u_cpu.rf_ram.memory\[105\]\[0\] u_cpu.rf_ram.memory\[106\]\[0\]
+ u_cpu.rf_ram.memory\[107\]\[0\] _01555_ _01531_ _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_99_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07916__A1 _03502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06719__A2 _02988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09814_ _00208_ io_in[4] u_cpu.rf_ram.memory\[41\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05078__S1 _01525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07392__A2 _03375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09745_ _00139_ io_in[4] u_cpu.rf_ram.memory\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09669__A1 _04636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06957_ _03104_ _03127_ _03130_ _00407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05908_ _02440_ _00045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09676_ u_cpu.rf_ram.memory\[23\]\[1\] _04832_ _04834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06888_ _02754_ _02768_ _03088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07144__A2 _03227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08341__A1 _03901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08627_ _02467_ u_arbiter.i_wb_cpu_rdt\[18\] _04216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05839_ _02391_ _02394_ _02398_ _02399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08892__A2 _04371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05250__S1 _01525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04902__A1 _01487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08558_ _03903_ _04153_ _04154_ _04155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_74_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07509_ _03316_ _03435_ _03440_ _00649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09772__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08489_ _04091_ _04092_ _00978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10520_ _00893_ io_in[4] u_cpu.rf_ram.memory\[115\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09099__S _02910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05002__S1 _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10451_ _00824_ io_in[4] u_cpu.rf_ram.memory\[34\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06407__A1 _02782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08947__A3 _04031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10382_ _00755_ io_in[4] u_cpu.rf_ram.memory\[38\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06958__A2 _03127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07855__B _01441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11105__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05630__A2 _02179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07907__A1 _02619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11003_ _01372_ io_in[4] u_cpu.rf_ram.memory\[26\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05069__S1 _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07383__A2 _03365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08580__B2 _04008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08332__A1 _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07135__A2 _03227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08883__A2 _04361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05241__S1 _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05697__A2 _02273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08635__A2 _02416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05449__A2 _02028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10718_ _01088_ io_in[4] u_cpu.rf_ram.memory\[109\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10649_ _01022_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08399__A1 _04009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09060__A2 _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06949__A2 _03117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07071__A1 _03110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05621__A2 _02198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07860_ _02285_ _02309_ _03639_ _03641_ _03643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07374__A2 _03365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06811_ _02657_ _03039_ _03045_ _00346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08571__B2 _04019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05385__A1 _01490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07791_ _03508_ _03593_ _03600_ _00771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08596__B _04031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09530_ u_cpu.rf_ram.memory\[27\]\[0\] _04752_ _04753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06742_ _02897_ _02998_ _03006_ _00316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05480__S1 _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10622__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08323__A1 _03936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07126__A2 _03217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09461_ u_cpu.rf_ram.memory\[87\]\[4\] _04701_ _04706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06673_ _02881_ _02967_ _02968_ _00285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09795__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08874__A2 _04361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06885__A1 _02895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08412_ u_arbiter.i_wb_cpu_rdt\[22\] u_arbiter.i_wb_cpu_rdt\[6\] _02466_ _04030_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05624_ u_cpu.rf_ram.memory\[52\]\[7\] u_cpu.rf_ram.memory\[53\]\[7\] u_cpu.rf_ram.memory\[54\]\[7\]
+ u_cpu.rf_ram.memory\[55\]\[7\] _01572_ _01573_ _02202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09392_ _04634_ _04661_ _04667_ _01306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05232__S1 _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08343_ _02313_ _03956_ _03958_ _03959_ _03968_ _00956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_51_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10772__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05555_ _01566_ _02133_ _01558_ _02134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08626__A2 _03910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06637__A1 _02885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08274_ _02465_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\] _03902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05486_ _01617_ _02065_ _01519_ _02066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06101__A3 _02585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07225_ _03102_ _03277_ _03279_ _00526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10002__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11128__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05860__A2 _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07156_ u_cpu.rf_ram.memory\[52\]\[3\] _03237_ _03241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05179__C _01560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06107_ _02586_ _02593_ _02596_ _00022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07087_ _03108_ _03197_ _03202_ _00465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06038_ _02538_ _02529_ _02528_ _02521_ _02539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__10152__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08562__A1 _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07365__A2 _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07989_ u_cpu.rf_ram.memory\[121\]\[0\] _03720_ _03721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09728_ _00122_ io_in[4] u_cpu.rf_ram.memory\[18\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08314__A1 _03940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07117__A2 _03217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09659_ _04626_ _04822_ _04824_ _01416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_76_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08865__A2 _04351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05223__S1 _01622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08726__S _02335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08617__A2 _03906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09290__A2 _04603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10503_ _00876_ io_in[4] u_cpu.rf_ram.memory\[112\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10434_ _00807_ io_in[4] u_cpu.rf_ram.memory\[92\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05851__A2 _02402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09042__A2 _04463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07053__A1 _03110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10365_ _00012_ io_in[4] u_cpu.rf_ram_if.rdata0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05603__A2 _02180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10296_ _00682_ io_in[4] u_cpu.rf_ram.memory\[130\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10645__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08553__A1 _03925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07356__A2 _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07108__A2 _03207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05119__A1 _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10795__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08856__A2 _04351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06867__A1 _02895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05214__S1 _01594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08608__A2 _04165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10025__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06619__A1 _02885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05340_ u_cpu.rf_ram.memory\[0\]\[4\] u_cpu.rf_ram.memory\[1\]\[4\] u_cpu.rf_ram.memory\[2\]\[4\]
+ u_cpu.rf_ram.memory\[3\]\[4\] _01530_ _01532_ _01921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__04963__I _01504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09281__A2 _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05271_ _01566_ _01852_ _01480_ _01853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_31_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07010_ u_cpu.rf_ram.memory\[19\]\[2\] _03157_ _03160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10175__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09033__A2 _04463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07595__A2 _03485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08170__I _03829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08961_ _03965_ _03962_ _04420_ _04421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_142_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07912_ _03498_ _03672_ _03674_ _00819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08892_ u_cpu.rf_ram.memory\[2\]\[0\] _04371_ _04372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07347__A2 _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07843_ u_cpu.rf_ram.memory\[90\]\[4\] _03626_ _03631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_04986_ _01463_ _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07774_ u_cpu.rf_ram.memory\[37\]\[7\] _03583_ _03591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09513_ _04739_ _04720_ _04740_ _01354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06725_ _02768_ _02803_ _02997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09444_ _04632_ _04691_ _04696_ _01329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06656_ _02885_ _02956_ _02958_ _00278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05905__I0 u_arbiter.i_wb_cpu_rdt\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05607_ _01528_ _02184_ _02185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05530__A1 _01463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06587_ u_cpu.cpu.state.genblk1.misalign_trap_sync_r u_cpu.cpu.state.stage_two_req
+ _02911_ _02912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09375_ u_cpu.rf_ram.memory\[10\]\[6\] _04651_ _04658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__04964__S0 _01495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08326_ _03897_ _03952_ _03953_ _00954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05538_ u_cpu.rf_ram.memory\[48\]\[6\] u_cpu.rf_ram.memory\[49\]\[6\] u_cpu.rf_ram.memory\[50\]\[6\]
+ u_cpu.rf_ram.memory\[51\]\[6\] _01576_ _01577_ _02117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_71_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09272__A2 _04593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10518__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08257_ _03699_ _03885_ _03889_ _00949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05469_ _01602_ _02048_ _02049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07208_ u_cpu.rf_ram.memory\[142\]\[2\] _03267_ _03270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05833__A2 _02392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08188_ _03844_ _03845_ _00924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09810__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09024__A2 _04453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07035__A1 _02657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07139_ _03106_ _03227_ _03231_ _00488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08232__B1 _03808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05046__B1 _01628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10668__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07586__A2 _03475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10150_ _00536_ io_in[4] u_cpu.rf_ram.memory\[140\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09960__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10081_ _00475_ io_in[4] u_cpu.rf_ram.memory\[55\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07338__A2 _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08535__A1 _03966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05653__B _01600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05444__S1 _01594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08838__A2 _04327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10983_ _01352_ io_in[4] u_cpu.cpu.genblk3.csr.mcause3_0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10048__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06849__A1 _02895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07510__A2 _03435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05521__A1 _01513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10198__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09263__A2 _02825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05824__A2 _01467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09015__A2 _04453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05380__S0 _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10417_ _00790_ io_in[4] u_cpu.rf_ram.memory\[90\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08223__B1 _03829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07577__A2 _03475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10348_ _00734_ io_in[4] u_cpu.rf_ram.memory\[124\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10279_ _00665_ io_in[4] u_cpu.rf_ram.memory\[132\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07329__A2 _03335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04958__I _01463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05435__S1 _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06510_ _02683_ _02861_ _02864_ _00226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07490_ u_cpu.rf_ram.memory\[135\]\[4\] _03425_ _03430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07501__A2 _03435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06441_ _02691_ _02816_ _02823_ _00198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05512__A1 _01506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09160_ _04438_ _04533_ _04535_ _01206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06372_ u_cpu.rf_ram.memory\[42\]\[0\] _02784_ _02785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09833__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09254__A2 _04583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08111_ u_cpu.rf_ram.memory\[116\]\[7\] _03780_ _03788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05323_ _01465_ _01904_ _01905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09091_ u_arbiter.i_wb_cpu_rdt\[27\] _04485_ _04497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07265__A1 _02647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08042_ _03749_ _03750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05254_ u_cpu.rf_ram.memory\[8\]\[3\] u_cpu.rf_ram.memory\[9\]\[3\] u_cpu.rf_ram.memory\[10\]\[3\]
+ u_cpu.rf_ram.memory\[11\]\[3\] _01523_ _01525_ _01836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10810__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05815__A2 _02274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05371__S0 _01529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07017__A1 _03110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09983__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08214__B1 _03829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05185_ _01571_ _01767_ _01768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08765__A1 _03691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07568__A2 _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09993_ _00387_ io_in[4] u_cpu.rf_ram.memory\[64\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10960__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06240__A2 _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08944_ _03945_ _03988_ _04188_ _04406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05674__S1 _01525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08875_ _02632_ _04361_ _04362_ _01094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09190__A1 _04450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07826_ _03504_ _03616_ _03621_ _00785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05426__S1 _01525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07740__A2 _03037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04969_ _01463_ _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05751__A1 _01445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07757_ _03510_ _03573_ _03581_ _00756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_77_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06708_ _02987_ _02988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07688_ u_cpu.rf_ram.memory\[125\]\[0\] _03543_ _03544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09427_ u_cpu.rf_ram.memory\[86\]\[5\] _04681_ _04687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10340__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06639_ _02887_ _02945_ _02948_ _00271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05503__A1 _02073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09358_ _04636_ _04641_ _04648_ _01291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09245__A2 _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08309_ _02466_ _02411_ _03937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06059__A2 _02397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07256__A1 _02731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09289_ u_cpu.rf_ram.memory\[108\]\[3\] _04603_ _04607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10490__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05362__S0 _01576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08205__B1 _03833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08756__A1 _02355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07559__A2 _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10202_ _00588_ io_in[4] u_cpu.rf_ram.memory\[143\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05114__S0 _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10133_ _00519_ io_in[4] u_cpu.rf_ram.memory\[142\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06231__A2 _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05665__S1 _01500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08508__A1 _03940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10064_ _00458_ io_in[4] u_cpu.rf_ram.memory\[57\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05990__A1 _02499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09706__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05383__B _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05417__S1 _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07731__A2 _03563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05742__A1 _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10966_ _01335_ io_in[4] u_cpu.rf_ram.memory\[87\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09856__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09484__A2 _04711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07495__A1 _03320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06298__A2 _02733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10897_ _01266_ io_in[4] u_cpu.rf_ram.memory\[108\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10833__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09236__A2 _04573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07247__A1 _03106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08295__I0 u_arbiter.i_wb_cpu_rdt\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05353__S0 _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10983__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06470__A2 _02840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05105__S0 _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06222__A2 _02679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05025__A3 _01609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05656__S1 _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10213__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06990_ u_cpu.rf_ram.memory\[60\]\[1\] _03147_ _03149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05941_ _02460_ _02461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09172__A1 _04450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08660_ _03699_ _04237_ _04241_ _01000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05872_ u_arbiter.i_wb_cpu_rdt\[7\] u_arbiter.i_wb_cpu_dbus_dat\[4\] _02418_ _02422_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_27_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05408__S1 _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07722__A2 _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07611_ _02636_ _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_93_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10363__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05733__A1 _01445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08591_ _03947_ _03904_ _04182_ _03955_ _04183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_53_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07542_ u_cpu.rf_ram.memory\[132\]\[3\] _03455_ _03459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09475__A2 _04711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07473_ _03316_ _03415_ _03420_ _00633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06289__A2 _02733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05740__C u_cpu.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09212_ _04434_ _04563_ _04564_ _01229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06424_ _02693_ _02805_ _02813_ _00191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09227__A2 _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07238__A1 _02814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09143_ u_cpu.rf_ram.memory\[103\]\[2\] _04523_ _04526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06355_ _02683_ _02770_ _02773_ _00162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05306_ _01881_ _01883_ _01885_ _01887_ _01486_ _01888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__07789__A2 _03593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09074_ _04488_ _01167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06286_ u_cpu.cpu.immdec.imm11_7\[4\] _02622_ _02730_ _02731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__05344__S0 _01530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08025_ u_cpu.rf_ram.memory\[11\]\[0\] _03740_ _03741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05237_ _01638_ _01819_ _01482_ _01820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06461__A2 _02829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05168_ u_cpu.rf_ram.memory\[12\]\[2\] u_cpu.rf_ram.memory\[13\]\[2\] u_cpu.rf_ram.memory\[14\]\[2\]
+ u_cpu.rf_ram.memory\[15\]\[2\] _01530_ _01532_ _01751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_103_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09729__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06213__A2 _02679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09976_ _00370_ io_in[4] u_cpu.rf_ram.memory\[66\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05099_ _01505_ _01682_ _01579_ _01683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07961__A2 _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08927_ _03955_ _04390_ _04391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10706__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08858_ u_cpu.rf_ram.memory\[109\]\[1\] _04351_ _04353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09879__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07713__A2 _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07809_ _02395_ _02259_ _03610_ _03612_ _00777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_29_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05724__A1 _02289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08789_ _04314_ _01056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__05724__B2 u_cpu.cpu.genblk3.csr.mstatus_mie vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10820_ _01189_ io_in[4] u_cpu.rf_ram.memory\[102\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10856__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09466__A2 _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07477__A1 _03320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10751_ _01120_ io_in[4] u_cpu.cpu.immdec.imm11_7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09218__A2 _04563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10682_ _00024_ io_in[4] u_cpu.cpu.ctrl.pc_plus_offset_cy_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08734__S _02335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07229__A1 _03106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08277__I0 u_arbiter.i_wb_cpu_rdt\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05335__S0 _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06452__A2 _02829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10236__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06204__A2 _02679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07401__A1 _03316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11165_ io_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_122_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07952__A2 _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10116_ _00510_ io_in[4] u_cpu.rf_ram.memory\[15\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11096_ _00094_ io_in[0] u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10386__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05963__A1 _02463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09154__A1 _04450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10047_ _00441_ io_in[4] u_cpu.rf_ram.memory\[5\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07704__A2 _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08901__A1 _02652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09457__A2 _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05560__C _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10949_ _01318_ io_in[4] u_cpu.rf_ram.memory\[86\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09209__A2 _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06140__A1 u_cpu.cpu.immdec.imm11_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11011__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06691__A2 _02978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08968__A1 _03691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06140_ u_cpu.cpu.immdec.imm11_7\[3\] _02620_ _02624_ _02625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_118_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04971__I _01498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06443__A2 _02816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06071_ u_scanchain_local.module_data_in\[64\] _02566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07640__A1 u_cpu.rf_ram.memory\[128\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05022_ _01518_ _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_126_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10729__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08196__A2 _03822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09830_ _00224_ io_in[4] u_cpu.rf_ram.memory\[48\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05403__B1 _01981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09761_ _00155_ io_in[4] u_cpu.rf_ram.memory\[80\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05954__A1 _02456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06973_ _03102_ _03137_ _03139_ _00414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08712_ u_arbiter.i_wb_cpu_dbus_adr\[13\] u_arbiter.i_wb_cpu_dbus_adr\[14\] _04257_
+ _04269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05924_ u_scanchain_local.module_data_in\[34\] u_arbiter.i_wb_cpu_dbus_dat\[29\]
+ _02431_ _02449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10879__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09692_ _04309_ _04841_ _04842_ _01431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_55_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08643_ u_arbiter.i_wb_cpu_rdt\[31\] u_arbiter.i_wb_cpu_rdt\[15\] _02467_ _04230_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_27_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05855_ u_arbiter.i_wb_cpu_rdt\[1\] _02411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05706__A1 _01441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08574_ _04167_ _04165_ _04168_ _03993_ _00987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_82_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09448__A2 _04691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05786_ _02359_ u_cpu.cpu.ctrl.i_iscomp _02360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10109__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07525_ _03314_ _03445_ _03449_ _00656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07459__A1 _03320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08120__A2 _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06131__A1 _01494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07456_ u_cpu.rf_ram.memory\[49\]\[5\] _03405_ _03411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06407_ _02782_ _02803_ _02804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06682__A2 _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10259__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07387_ _02662_ _03365_ _03372_ _00595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_109_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08959__A1 _03901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09126_ _04440_ _04513_ _04516_ _01191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06338_ u_cpu.rf_ram.memory\[80\]\[5\] _02756_ _02762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09620__A2 _04802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05198__B _01558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06269_ u_cpu.rf_ram.memory\[20\]\[1\] _02719_ _02721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06434__A2 _02816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07631__A1 _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09057_ _04440_ _04476_ _04479_ _01159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08008_ _02632_ _03730_ _03731_ _00858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09384__A1 _04626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08187__A2 _03822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07934__A2 _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09959_ _00353_ io_in[4] u_cpu.rf_ram.memory\[68\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09136__A1 _04450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09687__A2 _04832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09439__A2 _04691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06370__A1 _02780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11034__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10803_ _01172_ io_in[4] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08111__A2 _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10734_ _01103_ io_in[4] u_cpu.rf_ram.memory\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06122__A1 _02303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05556__S0 _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06673__A2 _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07870__A1 _02395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10665_ _01038_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10596_ _00969_ io_in[4] u_cpu.rf_ram.memory\[114\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09611__A2 _04792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07622__A1 _03504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05228__A3 _01810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08178__A2 _03822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07925__A2 _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11148_ _00082_ io_in[0] u_scanchain_local.module_data_in\[60\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11079_ u_cpu.rf_ram_if.wdata1_r\[3\] io_in[4] u_cpu.rf_ram_if.wdata1_r\[2\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09678__A2 _04832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07689__A1 _03494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08350__A2 _03947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__04966__I _01495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05640_ u_cpu.rf_ram.memory\[124\]\[7\] u_cpu.rf_ram.memory\[125\]\[7\] u_cpu.rf_ram.memory\[126\]\[7\]
+ u_cpu.rf_ram.memory\[127\]\[7\] _01496_ _01594_ _02218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06361__A1 _02689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05571_ u_cpu.rf_ram.memory\[64\]\[6\] u_cpu.rf_ram.memory\[65\]\[6\] u_cpu.rf_ram.memory\[66\]\[6\]
+ u_cpu.rf_ram.memory\[67\]\[6\] _01522_ _01622_ _02150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08102__A2 _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07310_ u_cpu.rf_ram.memory\[73\]\[4\] _03325_ _03330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10401__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08290_ _03906_ _03917_ _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05547__S0 _01529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07241_ _03098_ _03287_ _03288_ _00533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06664__A2 _02956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07172_ u_cpu.rf_ram.memory\[9\]\[2\] _03247_ _03250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08173__I _03808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09602__A2 _04792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10551__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06123_ _02606_ _02303_ _02608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07613__A1 _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06416__A2 _02805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08810__B1 _04311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06054_ _02552_ _00083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_99_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05005_ _01512_ _01589_ _01590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08169__A2 _03822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09366__A1 _02637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07916__A2 _03672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09813_ _00207_ io_in[4] u_cpu.rf_ram.memory\[51\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05927__A1 _02403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09118__A1 _04450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09744_ _00138_ io_in[4] u_cpu.rf_ram.memory\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06956_ u_cpu.rf_ram.memory\[62\]\[2\] _03127_ _03130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09669__A2 _04822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05037__I _01499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11057__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05907_ u_arbiter.i_wb_cpu_rdt\[24\] u_arbiter.i_wb_cpu_dbus_dat\[21\] _02431_ _02440_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09675_ _04622_ _04832_ _04833_ _01423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06887_ _02897_ _03079_ _03087_ _00380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08341__A2 _03963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05481__B _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08626_ _03974_ _03910_ _04212_ _04214_ _04215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05838_ _02388_ _02397_ _02398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08557_ _03925_ _03948_ _03962_ _04154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_70_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09917__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05769_ u_cpu.cpu.alu.i_rs1 _02277_ _02344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__04902__A2 _01488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10081__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07508_ u_cpu.rf_ram.memory\[134\]\[4\] _03435_ _03440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08488_ u_cpu.cpu.immdec.imm24_20\[4\] _04069_ _04070_ u_cpu.cpu.immdec.imm30_25\[0\]
+ _04088_ _04009_ _04092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__05538__S0 _01576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07852__A1 u_cpu.cpu.state.genblk1.misalign_trap_sync_r vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07439_ _03318_ _03395_ _03401_ _00618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06655__A2 _02956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10450_ _00823_ io_in[4] u_cpu.rf_ram.memory\[34\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09109_ u_cpu.rf_ram.memory\[101\]\[3\] _04503_ _04507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06407__A2 _02803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10381_ _00754_ io_in[4] u_cpu.rf_ram.memory\[38\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07080__A2 _03197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05091__B2 _01674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05630__A3 _02188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11002_ _01371_ io_in[4] u_cpu.rf_ram.memory\[26\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07907__A2 _02782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05375__C _01560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05918__A1 u_arbiter.i_wb_cpu_rdt\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08580__A2 _04165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08332__A2 u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10424__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06343__A1 _02693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06894__A2 _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05529__S0 _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10574__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10717_ _01087_ io_in[4] u_cpu.rf_ram.memory\[109\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06646__A2 _02945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10648_ _01021_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08399__A2 _04010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08643__I0 u_arbiter.i_wb_cpu_rdt\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10579_ _00952_ io_in[4] u_cpu.rf_ram.memory\[113\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07071__A2 _03187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09348__A1 _04626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08020__A1 _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06810_ u_cpu.rf_ram.memory\[6\]\[5\] _03039_ _03045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08571__A2 _04165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07790_ u_cpu.rf_ram.memory\[36\]\[6\] _03593_ _03600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05385__A2 _01956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08596__C _04051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06741_ u_cpu.rf_ram.memory\[77\]\[7\] _02998_ _03006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08323__A2 _03950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09460_ _04630_ _04701_ _04705_ _01336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06672_ u_cpu.rf_ram.memory\[119\]\[0\] _02967_ _02968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08411_ _01448_ _03956_ _04029_ _00963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05623_ _01548_ _02200_ _01480_ _02201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09391_ u_cpu.rf_ram.memory\[85\]\[5\] _04661_ _04667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06885__A2 _03079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10917__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08342_ _03960_ _03961_ _03967_ _03968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_71_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05554_ u_cpu.rf_ram.memory\[120\]\[6\] u_cpu.rf_ram.memory\[121\]\[6\] u_cpu.rf_ram.memory\[122\]\[6\]
+ u_cpu.rf_ram.memory\[123\]\[6\] _01598_ _01556_ _02133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_32_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06637__A2 _02945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08273_ _03900_ _03901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05485_ u_cpu.rf_ram.memory\[68\]\[5\] u_cpu.rf_ram.memory\[69\]\[5\] u_cpu.rf_ram.memory\[70\]\[5\]
+ u_cpu.rf_ram.memory\[71\]\[5\] _01507_ _01605_ _02065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_137_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07224_ u_cpu.rf_ram.memory\[141\]\[1\] _03277_ _03279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09587__A1 _04626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07155_ _03104_ _03237_ _03240_ _00495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06106_ _02594_ _02595_ _02596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07086_ u_cpu.rf_ram.memory\[56\]\[4\] _03197_ _03202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07062__A2 _03187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09339__A1 _04636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06037_ u_cpu.cpu.ctrl.o_ibus_adr\[20\] _02538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_133_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08562__A2 _03912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10447__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07988_ _03719_ _03720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06573__A1 _02642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09727_ _00121_ io_in[4] u_cpu.rf_ram.memory\[18\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06939_ _03104_ _03117_ _03120_ _00399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08314__A2 _03941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09658_ u_cpu.rf_ram.memory\[89\]\[1\] _04822_ _04824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10597__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08609_ _04165_ _04197_ _04198_ _04199_ _00991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__06876__A2 _03079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09589_ _04628_ _04782_ _04785_ _01385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04887__A1 u_cpu.cpu.immdec.imm19_12_20\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06628__A2 _02935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10502_ _00875_ io_in[4] u_cpu.rf_ram.memory\[112\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08742__S _02335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10433_ _00806_ io_in[4] u_cpu.rf_ram.memory\[92\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07053__A2 _03177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10364_ _00011_ io_in[4] u_cpu.rf_ram_if.rdata0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05064__A1 _01473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06800__A2 _03039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10295_ _00681_ io_in[4] u_cpu.rf_ram.memory\[130\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08002__A1 _03705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08553__A2 _03974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05206__I3 u_cpu.rf_ram.memory\[119\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08305__A2 _03932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06316__A1 _02647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06867__A2 _03069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07620__I _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05390__I2 u_cpu.rf_ram.memory\[82\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06619__A2 _02935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05270_ u_cpu.rf_ram.memory\[56\]\[3\] u_cpu.rf_ram.memory\[57\]\[3\] u_cpu.rf_ram.memory\[58\]\[3\]
+ u_cpu.rf_ram.memory\[59\]\[3\] _01567_ _01568_ _01852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_18_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07292__A2 _03308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09569__A1 _04626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07044__A2 _03177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05055__A1 _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08792__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08960_ _04024_ _04419_ _03948_ _04031_ _04420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_130_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07911_ u_cpu.rf_ram.memory\[34\]\[1\] _03672_ _03674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08891_ _04370_ _04371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09762__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07842_ _03502_ _03626_ _03630_ _00792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08400__B _04019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07773_ _03508_ _03583_ _03590_ _00763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_04985_ _01566_ _01569_ _01480_ _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_72_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09512_ u_cpu.cpu.genblk3.csr.mstatus_mie _04720_ _04740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_65_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06724_ _02897_ _02988_ _02996_ _00308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06307__A1 _02731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09443_ u_cpu.rf_ram.memory\[111\]\[4\] _04691_ _04696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06858__A2 _03069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06655_ u_cpu.rf_ram.memory\[40\]\[1\] _02956_ _02958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05606_ u_cpu.rf_ram.memory\[8\]\[7\] u_cpu.rf_ram.memory\[9\]\[7\] u_cpu.rf_ram.memory\[10\]\[7\]
+ u_cpu.rf_ram.memory\[11\]\[7\] _01497_ _01501_ _02184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_12_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09374_ _02657_ _04651_ _04657_ _01298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_40_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06586_ _02909_ u_arbiter.i_wb_cpu_ibus_adr\[1\] _02910_ _02911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_71_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04964__S1 _01499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08325_ _02265_ _03897_ _03953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07807__A1 _02395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05537_ _01571_ _02115_ _02116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08256_ u_cpu.rf_ram.memory\[113\]\[3\] _03885_ _03889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07283__A2 _03308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05468_ u_cpu.rf_ram.memory\[112\]\[5\] u_cpu.rf_ram.memory\[113\]\[5\] u_cpu.rf_ram.memory\[114\]\[5\]
+ u_cpu.rf_ram.memory\[115\]\[5\] _01572_ _01573_ _02048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08480__A1 u_cpu.cpu.immdec.imm24_20\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05050__I _01622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07207_ _03102_ _03267_ _03269_ _00518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08187_ u_arbiter.i_wb_cpu_rdt\[10\] _03822_ _03833_ u_arbiter.i_wb_cpu_dbus_dat\[11\]
+ _03845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_119_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05399_ u_cpu.rf_ram.memory\[72\]\[4\] u_cpu.rf_ram.memory\[73\]\[4\] u_cpu.rf_ram.memory\[74\]\[4\]
+ u_cpu.rf_ram.memory\[75\]\[4\] _01562_ _01622_ _01980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_119_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08232__A1 u_arbiter.i_wb_cpu_rdt\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07035__A2 _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07138_ u_cpu.rf_ram.memory\[53\]\[3\] _03227_ _03231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07069_ _03108_ _03187_ _03192_ _00457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06794__A1 _02895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10080_ _00474_ io_in[4] u_cpu.rf_ram.memory\[55\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08299__A1 _02464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10982_ _01351_ io_in[4] u_cpu.cpu.genblk3.csr.mcause3_0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06849__A2 _03059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09099__I0 u_arbiter.i_wb_cpu_rdt\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05521__A2 _02099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06077__A3 _02562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05380__S1 _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10612__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10416_ _00789_ io_in[4] u_cpu.rf_ram.memory\[90\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07026__A2 _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08223__A1 u_arbiter.i_wb_cpu_rdt\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09785__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08774__A2 _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10347_ _00733_ io_in[4] u_cpu.rf_ram.memory\[124\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10278_ _00664_ io_in[4] u_cpu.rf_ram.memory\[132\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10762__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06537__A1 _02691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11118__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05899__I0 u_arbiter.i_wb_cpu_rdt\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06440_ u_cpu.rf_ram.memory\[44\]\[6\] _02816_ _02823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10142__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06371_ _02783_ _02784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08110_ _03705_ _03780_ _03787_ _00904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05322_ u_cpu.rf_ram.memory\[136\]\[3\] u_cpu.rf_ram.memory\[137\]\[3\] u_cpu.rf_ram.memory\[138\]\[3\]
+ u_cpu.rf_ram.memory\[139\]\[3\] _01641_ _01642_ _01904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_119_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09090_ _04496_ _01175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07265__A2 _03297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08462__A1 _03955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08041_ _02754_ _02965_ _03749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05276__B2 _01857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05253_ _01528_ _01834_ _01534_ _01835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_70_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10292__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05371__S1 _01500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07017__A2 _03157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08214__A1 u_arbiter.i_wb_cpu_rdt\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05184_ u_cpu.rf_ram.memory\[52\]\[2\] u_cpu.rf_ram.memory\[53\]\[2\] u_cpu.rf_ram.memory\[54\]\[2\]
+ u_cpu.rf_ram.memory\[55\]\[2\] _01572_ _01573_ _01767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_143_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08765__A2 _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09992_ _00386_ io_in[4] u_cpu.rf_ram.memory\[64\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06776__A1 _02895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08943_ _03924_ _03977_ _03985_ _04405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_9_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08874_ u_cpu.rf_ram.memory\[3\]\[0\] _04361_ _04362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09190__A2 _04543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07825_ u_cpu.rf_ram.memory\[91\]\[4\] _03616_ _03621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__04929__I2 u_cpu.rf_ram.memory\[22\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07756_ u_cpu.rf_ram.memory\[38\]\[7\] _03573_ _03581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04968_ _01505_ _01552_ _01553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05751__A2 u_arbiter.i_wb_cpu_dbus_we vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06707_ _02849_ _02976_ _02987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07687_ _03542_ _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04899_ _01485_ _01486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_13_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09426_ _04632_ _04681_ _04686_ _01321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06638_ u_cpu.rf_ram.memory\[17\]\[2\] _02945_ _02948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06700__A1 _02891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05503__A2 _02082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09357_ u_cpu.rf_ram.memory\[59\]\[6\] _04641_ _04648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06569_ _02632_ _02900_ _02901_ _00248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_139_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10635__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08308_ _03933_ _03935_ _03936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07256__A2 _02803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09288_ _04440_ _04603_ _04606_ _01263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05267__A1 _01842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08239_ u_arbiter.i_wb_cpu_dbus_dat\[28\] _03808_ _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05362__S1 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07008__A2 _03157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08205__A1 u_arbiter.i_wb_cpu_rdt\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05648__C _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10785__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05019__A1 _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10201_ _00587_ io_in[4] u_cpu.rf_ram.memory\[143\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08756__A2 _04293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05114__S1 _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10132_ _00518_ io_in[4] u_cpu.rf_ram.memory\[142\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08508__A2 _03963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10015__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10063_ _00457_ io_in[4] u_cpu.rf_ram.memory\[57\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09181__A2 _04543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10165__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10965_ _01334_ io_in[4] u_cpu.rf_ram.memory\[87\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08141__B1 _03808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07495__A2 _03425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10896_ _01265_ io_in[4] u_cpu.rf_ram.memory\[108\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08444__A1 _04000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07247__A2 _03287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08995__A2 _04436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05839__B _02398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05353__S1 _01531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05105__S1 _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06758__A1 _02895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04969__I _01463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05574__B _01519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05940_ _02396_ u_cpu.cpu.state.ibus_cyc _02460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_67_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09172__A2 _04533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10508__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05871_ _02421_ _00095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_61_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07183__A1 _02667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07610_ _03494_ _03496_ _03497_ _00693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08590_ _03965_ _04175_ _04176_ _04181_ _04182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09800__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05733__A2 _02303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11090__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07541_ _03312_ _03455_ _03458_ _00663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10658__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07486__A2 _03425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07472_ u_cpu.rf_ram.memory\[136\]\[4\] _03415_ _03420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09211_ u_cpu.rf_ram.memory\[105\]\[0\] _04563_ _04564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05497__A1 _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06423_ u_cpu.rf_ram.memory\[45\]\[7\] _02805_ _02813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09950__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09142_ _04438_ _04523_ _04525_ _01198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06354_ u_cpu.rf_ram.memory\[78\]\[2\] _02770_ _02773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07238__A2 _02976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05305_ _01617_ _01886_ _01607_ _01887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08986__A2 _04436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09073_ u_arbiter.i_wb_cpu_rdt\[18\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[2\]
+ _04485_ _04488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06285_ _02728_ _02608_ _02729_ _02730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06997__A1 _03108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05344__S1 _01532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08024_ _03739_ _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05236_ u_cpu.rf_ram.memory\[132\]\[2\] u_cpu.rf_ram.memory\[133\]\[2\] u_cpu.rf_ram.memory\[134\]\[2\]
+ u_cpu.rf_ram.memory\[135\]\[2\] _01641_ _01642_ _01819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08199__B1 _03833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10038__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05167_ _01528_ _01749_ _01750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05098_ u_cpu.rf_ram.memory\[48\]\[1\] u_cpu.rf_ram.memory\[49\]\[1\] u_cpu.rf_ram.memory\[50\]\[1\]
+ u_cpu.rf_ram.memory\[51\]\[1\] _01576_ _01577_ _01682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07410__A2 _03385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09975_ _00369_ io_in[4] u_cpu.rf_ram.memory\[66\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08926_ _02392_ _02604_ _04390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_131_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09163__A2 _04533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10188__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08857_ _03691_ _04351_ _04352_ _01086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_18_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08910__A2 _04381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07808_ u_cpu.cpu.state.o_cnt_r\[3\] _03611_ _03612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08788_ u_cpu.cpu.ctrl.o_ibus_adr\[2\] _04309_ _04311_ u_cpu.cpu.ctrl.o_ibus_adr\[3\]
+ _04314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05724__A2 _02276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07739_ _03510_ _03563_ _03571_ _00748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10750_ _01119_ io_in[4] u_cpu.cpu.immdec.imm11_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08674__A1 _03695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07477__A2 _03415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05488__A1 _01621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09409_ u_cpu.rf_ram.memory\[110\]\[5\] _04671_ _04677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10681_ _01053_ io_in[4] u_cpu.rf_ram.memory\[30\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08426__A1 _03691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07229__A2 _03277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08977__A2 _04425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05335__S1 _01509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05660__A1 _01621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07401__A2 _03375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11164_ io_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_96_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10115_ _00509_ io_in[4] u_cpu.rf_ram.memory\[15\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11095_ _00093_ io_in[0] u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09823__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09154__A2 _04523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10046_ _00440_ io_in[4] u_cpu.rf_ram.memory\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07165__A1 _03114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08901__A2 _04371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09380__I _04660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10800__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05566__I2 u_cpu.rf_ram.memory\[82\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09973__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10948_ _01317_ io_in[4] u_cpu.rf_ram.memory\[86\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07468__A2 _03415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05479__A1 _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10950__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10879_ _01248_ io_in[4] u_cpu.rf_ram.memory\[107\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08417__A1 _03986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08968__A2 _04425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05569__B _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06979__A1 _03108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06070_ _02562_ _02564_ _02565_ _00086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07640__A2 _03513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05651__A1 _01464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05021_ u_cpu.rf_ram.memory\[116\]\[0\] u_cpu.rf_ram.memory\[117\]\[0\] u_cpu.rf_ram.memory\[118\]\[0\]
+ u_cpu.rf_ram.memory\[119\]\[0\] _01576_ _01605_ _01606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_144_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09393__A2 _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10330__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09760_ _00154_ io_in[4] u_cpu.rf_ram.memory\[80\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06972_ u_cpu.rf_ram.memory\[61\]\[1\] _03137_ _03139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08711_ _04268_ _01024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09145__A2 _04523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05923_ _02448_ _00053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09691_ u_cpu.cpu.state.ibus_cyc _04841_ _04842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_27_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08642_ _04165_ _04226_ _04228_ _04229_ _00994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_54_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10480__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05854_ _02410_ _00059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06903__A1 _02895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05706__A2 u_cpu.cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08573_ u_cpu.cpu.immdec.imm19_12_20\[2\] _03897_ _04165_ _04168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05785_ u_cpu.cpu.state.o_cnt_r\[1\] _02359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07524_ u_cpu.rf_ram.memory\[133\]\[3\] _03445_ _03449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07459__A2 _03405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08656__A1 _03695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05014__S0 _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07455_ _03316_ _03405_ _03410_ _00625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06406_ _02672_ _02765_ _02803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08408__A1 _03938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08408__B2 _03944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07386_ u_cpu.rf_ram.memory\[14\]\[6\] _03365_ _03372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_124_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09125_ u_cpu.rf_ram.memory\[102\]\[2\] _04513_ _04516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06337_ _02687_ _02756_ _02761_ _00156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09056_ u_cpu.rf_ram.memory\[28\]\[2\] _04476_ _04479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06268_ _02669_ _02719_ _02720_ _00128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07631__A2 _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08007_ u_cpu.rf_ram.memory\[8\]\[0\] _03730_ _03731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05219_ u_cpu.rf_ram.memory\[64\]\[2\] u_cpu.rf_ram.memory\[65\]\[2\] u_cpu.rf_ram.memory\[66\]\[2\]
+ u_cpu.rf_ram.memory\[67\]\[2\] _01522_ _01622_ _01802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_116_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06199_ u_cpu.cpu.immdec.imm11_7\[3\] u_cpu.cpu.immdec.imm11_7\[4\] _02620_ _02622_
+ _02676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_104_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09846__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09384__A2 _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07395__A1 _03310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09958_ _00352_ io_in[4] u_cpu.rf_ram.memory\[68\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10823__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09136__A2 _04513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08909_ _04380_ _04381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_106_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07147__A1 _03114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09889_ _00283_ io_in[4] u_cpu.rf_ram.memory\[40\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09996__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07698__A2 _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08895__A1 _02637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10973__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06370__A2 _02782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10802_ _01171_ io_in[4] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10733_ _01102_ io_in[4] u_cpu.rf_ram.memory\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05556__S1 _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10203__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10664_ _01037_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05389__B _01600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10595_ _00968_ io_in[4] u_cpu.rf_ram.memory\[114\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07622__A2 _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10353__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09375__A2 _04651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11147_ _00080_ io_in[0] u_scanchain_local.module_data_in\[59\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09127__A2 _04513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11078_ u_cpu.rf_ram_if.wdata1_r\[2\] io_in[4] u_cpu.rf_ram_if.wdata1_r\[1\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10029_ _00423_ io_in[4] u_cpu.rf_ram.memory\[60\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07689__A2 _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07623__I _02656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06361__A2 _02770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05570_ _02142_ _02144_ _02146_ _02148_ _01486_ _02149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_91_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08638__A1 _03922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09719__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05547__S1 _01500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04982__I _01494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07240_ u_cpu.rf_ram.memory\[140\]\[0\] _03287_ _03288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07171_ _02637_ _03247_ _03249_ _00502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09063__A1 _04446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09869__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06122_ _02303_ _01455_ _02607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__08390__S _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07613__A2 _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08810__B2 u_cpu.cpu.ctrl.o_ibus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06053_ _02389_ u_scanchain_local.module_data_in\[60\] _02551_ _02552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10846__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05004_ u_cpu.rf_ram.memory\[108\]\[0\] u_cpu.rf_ram.memory\[109\]\[0\] u_cpu.rf_ram.memory\[110\]\[0\]
+ u_cpu.rf_ram.memory\[111\]\[0\] _01551_ _01524_ _01589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09366__A2 _04651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07377__A1 _02637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09812_ _00206_ io_in[4] u_cpu.rf_ram.memory\[51\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09118__A2 _04503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05483__S0 _01522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09743_ _00137_ io_in[4] u_cpu.rf_ram.memory\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06955_ _03102_ _03127_ _03129_ _00406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07129__A1 _03114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10996__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05906_ _02439_ _00044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09674_ u_cpu.rf_ram.memory\[23\]\[0\] _04832_ _04833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06886_ u_cpu.rf_ram.memory\[65\]\[7\] _03079_ _03087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08877__A1 _02637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08625_ _03923_ _04052_ _04213_ _03915_ _04214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05837_ _02396_ u_cpu.cpu.state.ibus_cyc _02397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06352__A2 _02770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10226__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08629__A1 _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08556_ _03933_ _04000_ _03949_ _04153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05768_ _02305_ _02341_ _02342_ _02343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05053__I _01621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07507_ _03314_ _03435_ _03439_ _00648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08487_ _03966_ _04087_ _04089_ _04090_ _04091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_05699_ _02272_ _02274_ _02275_ _02276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05538__S1 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07438_ u_cpu.rf_ram.memory\[137\]\[5\] _03395_ _03401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07852__A2 _03611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10376__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05863__A1 u_arbiter.i_wb_cpu_dbus_dat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07369_ _03320_ _03355_ _03362_ _00587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09108_ _04440_ _04503_ _04506_ _01183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07604__A2 _03485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10380_ _00753_ io_in[4] u_cpu.rf_ram.memory\[38\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09039_ u_cpu.rf_ram.memory\[96\]\[5\] _04463_ _04469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09357__A2 _04641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11001_ _01370_ io_in[4] u_cpu.rf_ram.memory\[26\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05918__A2 _02403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09109__A2 _04503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05474__S0 _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11001__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06591__A2 _02914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06343__A2 _02756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11151__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10719__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05529__S1 _01531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10716_ _01086_ io_in[4] u_cpu.rf_ram.memory\[109\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07843__A2 _03626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09045__A1 u_cpu.cpu.bufreg.i_sh_signed vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10647_ _01020_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10869__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09596__A2 _04782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10578_ _00951_ io_in[4] u_cpu.rf_ram.memory\[113\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08643__I1 u_arbiter.i_wb_cpu_rdt\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05847__B _02388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09348__A2 _04641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07359__A1 _03310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08020__A2 _03730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06031__A1 _02388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05385__A3 _01965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06582__A2 _02900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06740_ _02895_ _02998_ _03005_ _00315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10249__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08859__A1 _03695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04977__I _01495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09520__A2 _01477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06671_ _02966_ _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_64_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07531__A1 _03320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06334__A2 _02756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08410_ _04009_ _04020_ _04028_ _03955_ _04029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_58_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05622_ u_cpu.rf_ram.memory\[56\]\[7\] u_cpu.rf_ram.memory\[57\]\[7\] u_cpu.rf_ram.memory\[58\]\[7\]
+ u_cpu.rf_ram.memory\[59\]\[7\] _01567_ _01568_ _02200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09390_ _04632_ _04661_ _04666_ _01305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10399__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08341_ _03901_ _03963_ _03966_ _03967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__04896__A2 _01438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05553_ _01543_ _02131_ _02132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09284__A1 _04434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08087__A2 _03770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__04926__B _01481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08272_ u_arbiter.i_wb_cpu_rdt\[0\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[0\]
+ _02465_ _03900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_60_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05484_ _01621_ _02063_ _02064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05845__A1 _02403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07223_ _03098_ _03277_ _03278_ _00525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09036__A1 _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09587__A2 _04782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07154_ u_cpu.rf_ram.memory\[52\]\[2\] _03237_ _03240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06105_ u_cpu.cpu.state.stage_two_req _02315_ _02595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07085_ _03106_ _03197_ _03201_ _00464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06270__A1 _02681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09339__A2 _04624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06036_ _02463_ _02536_ _02537_ _00079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11024__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08011__A2 _03730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07987_ _02838_ _02965_ _03719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06573__A2 _02900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09726_ _00120_ io_in[4] u_cpu.rf_ram.memory\[18\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06938_ u_cpu.rf_ram.memory\[63\]\[2\] _03117_ _03120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06869_ _02897_ _03069_ _03077_ _00372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09657_ _04622_ _04822_ _04823_ _01415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08608_ u_cpu.cpu.immdec.imm19_12_20\[5\] _04165_ _04199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09588_ u_cpu.rf_ram.memory\[24\]\[2\] _04782_ _04785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08295__S _02464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08539_ _03923_ _03935_ _03922_ _04137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__04887__A2 u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07825__A2 _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10501_ _00874_ io_in[4] u_cpu.rf_ram.memory\[112\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09027__A1 _02754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09578__A2 _04772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10432_ _00805_ io_in[4] u_cpu.rf_ram.memory\[92\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08786__B1 _04311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10363_ _00010_ io_in[4] u_cpu.rf_ram_if.rdata0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08250__A2 _03885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10294_ _00680_ io_in[4] u_cpu.rf_ram.memory\[130\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08002__A2 _03720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06564__A2 _02883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07761__A1 _03494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08269__I _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09502__A2 _02303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10541__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07513__A1 _03320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06316__A2 _02745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08069__A2 _03760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09266__A1 _04434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08313__I0 u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10691__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05827__A1 _01467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09018__A1 _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09569__A2 _04772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11047__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06252__A1 _02683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05055__A2 _01639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05296__C _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07910_ _03494_ _03672_ _03673_ _00818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09907__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10071__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08890_ _02619_ _02731_ _04370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_68_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06004__A1 _02463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07841_ u_cpu.rf_ram.memory\[90\]\[3\] _03626_ _03630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06555__A2 _02883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07772_ u_cpu.rf_ram.memory\[37\]\[6\] _03583_ _03590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04984_ u_cpu.rf_ram.memory\[56\]\[0\] u_cpu.rf_ram.memory\[57\]\[0\] u_cpu.rf_ram.memory\[58\]\[0\]
+ u_cpu.rf_ram.memory\[59\]\[0\] _01567_ _01568_ _01569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09511_ u_cpu.cpu.genblk3.csr.mstatus_mpie _04739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06723_ u_cpu.rf_ram.memory\[139\]\[7\] _02988_ _02996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06307__A2 _02743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09442_ _04630_ _04691_ _04695_ _01328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_92_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06654_ _02881_ _02956_ _02957_ _00277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05605_ _01528_ _02182_ _01534_ _02183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09373_ u_cpu.rf_ram.memory\[10\]\[5\] _04651_ _04657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06585_ u_arbiter.i_wb_cpu_ack _02461_ _02910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08304__I0 u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08324_ _03899_ _03912_ _03915_ _03931_ _03951_ _03952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_21_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05536_ u_cpu.rf_ram.memory\[52\]\[6\] u_cpu.rf_ram.memory\[53\]\[6\] u_cpu.rf_ram.memory\[54\]\[6\]
+ u_cpu.rf_ram.memory\[55\]\[6\] _01572_ _01573_ _02115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07807__A2 _02263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09009__A1 _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08255_ _03697_ _03885_ _03888_ _00948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05467_ _01566_ _02046_ _01600_ _02047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08480__A2 _04069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07206_ u_cpu.rf_ram.memory\[142\]\[1\] _03267_ _03269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08186_ u_arbiter.i_wb_cpu_dbus_dat\[10\] _03835_ _03844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05398_ _01617_ _01978_ _01519_ _01979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_4_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07137_ _03104_ _03227_ _03230_ _00487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08232__A2 _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10414__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07068_ u_cpu.rf_ram.memory\[57\]\[4\] _03187_ _03192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06794__A2 _03028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06019_ _02388_ _02522_ _02523_ _02524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_59_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10564__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06546__A2 _02883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07743__A1 _03494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06111__B _02599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09709_ _00103_ io_in[4] u_cpu.rf_ram.memory\[82\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10981_ _01350_ io_in[4] u_cpu.cpu.genblk3.csr.mcause3_0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09248__A1 _04434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09099__I1 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08456__C1 _03985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05809__A1 _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10415_ _00788_ io_in[4] u_cpu.rf_ram.memory\[91\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09420__A1 _04626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08223__A2 _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10094__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06234__A1 _02683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10346_ _00732_ io_in[4] u_cpu.rf_ram.memory\[125\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07982__A1 _03703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06785__A2 _03028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10907__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10277_ _00663_ io_in[4] u_cpu.rf_ram.memory\[132\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06537__A2 _02872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08931__B1 _03988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09487__A1 _02263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05860__B _02355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06370_ _02780_ _02782_ _02783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05321_ _01638_ _01902_ _01482_ _01903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08462__A2 _04068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10437__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06473__A1 _02683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08040_ _02667_ _03740_ _03748_ _00873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05276__A2 _01853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05252_ u_cpu.rf_ram.memory\[0\]\[3\] u_cpu.rf_ram.memory\[1\]\[3\] u_cpu.rf_ram.memory\[2\]\[3\]
+ u_cpu.rf_ram.memory\[3\]\[3\] _01530_ _01532_ _01834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_134_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08214__A2 _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05183_ _01566_ _01765_ _01480_ _01766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06225__A1 _02693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05659__S0 _01522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10587__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09991_ _00385_ io_in[4] u_cpu.rf_ram.memory\[64\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06776__A2 _03018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08942_ _03924_ _04403_ _04404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08411__B _04029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08873_ _04360_ _04361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07725__A1 _03494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06528__A2 _02872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07824_ _03502_ _03616_ _03620_ _00784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09478__A1 _04630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04967_ u_cpu.rf_ram.memory\[40\]\[0\] u_cpu.rf_ram.memory\[41\]\[0\] u_cpu.rf_ram.memory\[42\]\[0\]
+ u_cpu.rf_ram.memory\[43\]\[0\] _01551_ _01524_ _01552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_37_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07755_ _03508_ _03573_ _03580_ _00755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08525__I0 u_arbiter.i_wb_cpu_rdt\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06706_ _02897_ _02978_ _02986_ _00300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07686_ _02803_ _02965_ _03542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04898_ _01483_ _01484_ _01485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_44_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09425_ u_cpu.rf_ram.memory\[86\]\[4\] _04681_ _04686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06637_ _02885_ _02945_ _02947_ _00270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06700__A2 _02978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06568_ u_cpu.rf_ram.memory\[4\]\[0\] _02900_ _02901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09356_ _04634_ _04641_ _04647_ _01290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08307_ _02909_ u_arbiter.i_wb_cpu_rdt\[12\] _03934_ _03935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05519_ _01528_ _02097_ _02098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09287_ u_cpu.rf_ram.memory\[108\]\[2\] _04603_ _04606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06499_ u_cpu.rf_ram.memory\[43\]\[6\] _02851_ _02858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05267__A2 _01844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08238_ _03877_ _03878_ _00941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06464__A1 _02693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08169_ u_arbiter.i_wb_cpu_rdt\[5\] _03822_ _03832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09402__A1 _04626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08205__A2 _03822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06216__A1 _02687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10200_ _00586_ io_in[4] u_cpu.rf_ram.memory\[143\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06767__A2 _03018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10131_ _00517_ io_in[4] u_cpu.rf_ram.memory\[142\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10062_ _00456_ io_in[4] u_cpu.rf_ram.memory\[57\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06519__A2 _02861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07192__A2 _03257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09469__A1 _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04950__A1 _01528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10964_ _01333_ io_in[4] u_cpu.rf_ram.memory\[87\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08141__A1 u_arbiter.i_wb_cpu_rdt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08141__B2 u_arbiter.i_wb_cpu_dbus_dat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10895_ _01264_ io_in[4] u_cpu.rf_ram.memory\[108\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09641__A1 _04626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08444__A2 _04052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09752__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06207__A1 _02681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06758__A2 _03008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10329_ _00715_ io_in[4] u_cpu.rf_ram.memory\[127\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05966__B1 _02398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07626__I _02661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07707__A1 _03494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05870_ u_arbiter.i_wb_cpu_rdt\[6\] u_arbiter.i_wb_cpu_dbus_dat\[3\] _02418_ _02421_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07183__A2 _03247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05194__A1 _01548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06930__A2 _03100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07540_ u_cpu.rf_ram.memory\[132\]\[2\] _03455_ _03458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08132__A1 u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07471_ _03314_ _03415_ _03419_ _00632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08683__A2 _04247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09210_ _04562_ _04563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06422_ _02691_ _02805_ _02812_ _00190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05497__A2 _02076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06694__A1 _02885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09141_ u_cpu.rf_ram.memory\[103\]\[1\] _04523_ _04525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06353_ _02681_ _02770_ _02772_ _00161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08435__A2 _04041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08406__B _03938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05304_ u_cpu.rf_ram.memory\[84\]\[3\] u_cpu.rf_ram.memory\[85\]\[3\] u_cpu.rf_ram.memory\[86\]\[3\]
+ u_cpu.rf_ram.memory\[87\]\[3\] _01507_ _01605_ _01886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09072_ _04487_ _01166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06284_ u_cpu.cpu.immdec.imm11_7\[3\] _02608_ _02729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06997__A2 _03147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08023_ _02731_ _02849_ _03739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05235_ _01465_ _01817_ _01818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08199__A1 u_arbiter.i_wb_cpu_rdt\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05166_ u_cpu.rf_ram.memory\[8\]\[2\] u_cpu.rf_ram.memory\[9\]\[2\] u_cpu.rf_ram.memory\[10\]\[2\]
+ u_cpu.rf_ram.memory\[11\]\[2\] _01523_ _01525_ _01749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_115_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06749__A2 _03008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09974_ _00368_ io_in[4] u_cpu.rf_ram.memory\[66\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05957__B1 _02398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05097_ _01571_ _01680_ _01681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08925_ _03707_ _04381_ _04389_ _01117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08856_ u_cpu.rf_ram.memory\[109\]\[0\] _04351_ _04352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05056__I _01522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07174__A2 _03247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08371__A1 _02286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07807_ _02395_ _02263_ _03611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05185__A1 _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08787_ _04313_ _01055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_05999_ u_cpu.cpu.ctrl.o_ibus_adr\[13\] u_cpu.cpu.ctrl.o_ibus_adr\[12\] _02499_ _02508_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_55_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06921__A2 _03100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04895__I _01481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07738_ u_cpu.rf_ram.memory\[123\]\[7\] _03563_ _03571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10602__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07669_ _03532_ _03533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08674__A2 _04247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09775__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09408_ _04632_ _04671_ _04676_ _01313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06685__A1 _02895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10680_ _01052_ io_in[4] u_cpu.rf_ram.memory\[30\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09339_ _04636_ _04624_ _04637_ _01283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10752__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09623__A1 _04626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08426__A2 _04041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06437__A1 _02687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06988__A2 _03147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04999__A1 _01492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11108__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05660__A2 _02237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11163_ io_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_10114_ _00508_ io_in[4] u_cpu.rf_ram.memory\[9\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05394__C _01486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11094_ _00092_ io_in[0] u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10132__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10045_ _00439_ io_in[4] u_cpu.rf_ram.memory\[5\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08362__A1 _03974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07165__A2 _03237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05176__A1 _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06912__A2 _03100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10282__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10947_ _01316_ io_in[4] u_cpu.rf_ram.memory\[110\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08665__A2 _04237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05479__A2 _02058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06676__A1 u_cpu.rf_ram.memory\[119\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10878_ _01247_ io_in[4] u_cpu.rf_ram.memory\[107\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06979__A2 _03137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05100__B2 _01683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05020_ _01498_ _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05651__A2 _02228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07928__A1 _03494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05585__B _01482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06971_ _03098_ _03137_ _03138_ _00413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08710_ u_arbiter.i_wb_cpu_dbus_adr\[12\] u_arbiter.i_wb_cpu_dbus_adr\[13\] _04257_
+ _04268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05922_ u_arbiter.i_wb_cpu_rdt\[31\] u_arbiter.i_wb_cpu_dbus_dat\[28\] _02431_ _02448_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09690_ _03896_ _03611_ _04841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10625__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07156__A2 _03237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05853_ u_arbiter.i_wb_cpu_rdt\[0\] _02389_ _02409_ _02410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08641_ u_cpu.cpu.immdec.imm19_12_20\[8\] _04165_ _04229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05167__A1 _01528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09798__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06903__A2 _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08572_ u_cpu.cpu.immdec.imm19_12_20\[1\] _04167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05784_ _01442_ _02357_ _01444_ _02265_ _02358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07523_ _03312_ _03445_ _03448_ _00655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10775__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08656__A2 _04237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05014__S1 _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07454_ u_cpu.rf_ram.memory\[49\]\[4\] _03405_ _03410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09520__B _02303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06405_ _02693_ _02794_ _02802_ _00183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07385_ _02657_ _03365_ _03371_ _00594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10005__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09605__A1 _02681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09124_ _04438_ _04513_ _04515_ _01190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06336_ u_cpu.rf_ram.memory\[80\]\[4\] _02756_ _02761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09055_ _04438_ _04476_ _04478_ _01158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06267_ u_cpu.rf_ram.memory\[20\]\[0\] _02719_ _02720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05218_ _01794_ _01796_ _01798_ _01800_ _01486_ _01801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_08006_ _03729_ _03730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10155__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06198_ _02672_ _02674_ _02675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05149_ _01638_ _01732_ _01534_ _01733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07395__A2 _03375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08592__A1 u_cpu.cpu.immdec.imm19_12_20\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05245__I2 u_cpu.rf_ram.memory\[22\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09957_ _00351_ io_in[4] u_cpu.rf_ram.memory\[68\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08908_ _02626_ _02803_ _04380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09888_ _00282_ io_in[4] u_cpu.rf_ram.memory\[40\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08344__A1 _03901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07147__A2 _03227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05158__A1 _01513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08839_ _04340_ _01080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_57_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08895__A2 _04371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__04905__A1 _01465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10801_ _01170_ io_in[4] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06658__A1 _02887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10732_ _01101_ io_in[4] u_cpu.rf_ram.memory\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05330__A1 _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10663_ _01036_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10594_ _00967_ io_in[4] u_cpu.rf_ram.memory\[114\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07083__A1 _03104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11080__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10648__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07386__A2 _03365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11146_ _00079_ io_in[0] u_scanchain_local.module_data_in\[58\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09940__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11077_ u_cpu.rf_ram_if.wdata1_r\[1\] io_in[4] u_cpu.rf_ram_if.wdata1_r\[0\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08335__A1 _03914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07138__A2 _03227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10028_ _00422_ io_in[4] u_cpu.rf_ram.memory\[60\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05149__A1 _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10798__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08886__A2 _04361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06897__A1 _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10028__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06649__A1 _02897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07310__A2 _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05321__A1 _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07170_ u_cpu.rf_ram.memory\[9\]\[1\] _03247_ _03249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09063__A2 _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10178__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06121_ u_cpu.rf_ram_if.genblk1.wtrig0_r _02606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08810__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06052_ _02547_ _02549_ _02550_ _02388_ _02551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__06821__A1 _02885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05180__S0 _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05003_ _01548_ _01587_ _01579_ _01588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_67_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07377__A2 _03365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08574__B2 _03993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09811_ _00205_ io_in[4] u_cpu.rf_ram.memory\[51\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09742_ _00136_ io_in[4] u_cpu.rf_ram.memory\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05483__S1 _01622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06954_ u_cpu.rf_ram.memory\[62\]\[1\] _03127_ _03129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08326__A1 _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07129__A2 _03217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05905_ u_arbiter.i_wb_cpu_rdt\[23\] u_arbiter.i_wb_cpu_dbus_dat\[20\] _02431_ _02439_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09673_ _04831_ _04832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06885_ _02895_ _03079_ _03086_ _00379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08877__A2 _04361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06888__A1 _02754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08624_ _03918_ _03975_ _04013_ _04213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_54_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05836_ _02395_ _02396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_54_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08555_ _03935_ _03962_ _04151_ _04152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05767_ _02305_ _02317_ _02342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_78_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05560__A1 _02132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07506_ u_cpu.rf_ram.memory\[134\]\[3\] _03435_ _03439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08486_ _03914_ _03940_ _03938_ _04090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05698_ u_cpu.rf_ram_if.rdata1\[0\] _02272_ _02275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05312__A1 _01621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07437_ _03316_ _03395_ _03400_ _00617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05863__A2 _02389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06165__I _02646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09054__A2 _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07368_ u_cpu.rf_ram.memory\[143\]\[6\] _03355_ _03362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09813__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09107_ u_cpu.rf_ram.memory\[101\]\[2\] _04503_ _04506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07065__A1 _03104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06319_ u_cpu.rf_ram.memory\[7\]\[5\] _02745_ _02751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_136_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07299_ _03322_ _03308_ _03323_ _00556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09038_ _04444_ _04463_ _04468_ _01151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05171__S0 _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09963__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07368__A2 _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11000_ _01369_ io_in[4] u_cpu.rf_ram.memory\[26\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05379__A1 _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10940__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05474__S1 _01563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08868__A2 _04351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06879__A1 _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07540__A2 _03455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09293__A2 _04603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10320__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05303__A1 _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10715_ _01085_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10646_ _01019_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09045__A2 _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10577_ _00950_ io_in[4] u_cpu.rf_ram.memory\[113\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10470__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06803__A1 _02637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05162__S0 _01523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07359__A2 _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11129_ _00061_ io_in[0] u_scanchain_local.module_data_in\[41\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08859__A2 _04351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05790__A1 _01445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06670_ _02743_ _02965_ _02966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07531__A2 _03445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05621_ _01543_ _02198_ _02199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05542__A1 _01492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05552_ u_cpu.rf_ram.memory\[124\]\[6\] u_cpu.rf_ram.memory\[125\]\[6\] u_cpu.rf_ram.memory\[126\]\[6\]
+ u_cpu.rf_ram.memory\[127\]\[6\] _01496_ _01594_ _02131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08340_ _02911_ _03965_ _03966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09836__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09284__A2 _04603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08271_ _02465_ _02414_ _03898_ _03899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05483_ u_cpu.rf_ram.memory\[64\]\[5\] u_cpu.rf_ram.memory\[65\]\[5\] u_cpu.rf_ram.memory\[66\]\[5\]
+ u_cpu.rf_ram.memory\[67\]\[5\] _01522_ _01622_ _02063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_60_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05845__A2 u_cpu.cpu.genblk3.csr.i_mtip vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07222_ u_cpu.rf_ram.memory\[141\]\[0\] _03277_ _03278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10813__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09036__A2 _04463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07153_ _03102_ _03237_ _03239_ _00494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07047__A1 _03104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09986__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06104_ _02308_ _02312_ _02594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07598__A2 _03485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07084_ u_cpu.rf_ram.memory\[56\]\[3\] _03197_ _03201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05153__S0 _01497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10963__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06035_ _02402_ u_scanchain_local.module_data_in\[57\] _02478_ u_arbiter.i_wb_cpu_dbus_adr\[20\]
+ _02537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06270__A2 _02719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08547__A1 _02320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07986_ _03707_ _03710_ _03718_ _00849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07770__A2 _03583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09725_ _00119_ io_in[4] u_cpu.rf_ram.memory\[81\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06937_ _03102_ _03117_ _03119_ _00398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_41_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09656_ u_cpu.rf_ram.memory\[89\]\[0\] _04822_ _04823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06868_ u_cpu.rf_ram.memory\[66\]\[7\] _03069_ _03077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07522__A2 _03445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10343__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08607_ u_cpu.cpu.immdec.imm19_12_20\[6\] _03955_ _04198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_43_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05819_ _01467_ _02371_ _02383_ _00010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09587_ _04626_ _04782_ _04784_ _01384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__04967__S0 _01551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05533__A1 _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06799_ _03038_ _03039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08538_ u_arbiter.i_wb_cpu_rdt\[30\] u_arbiter.i_wb_cpu_rdt\[14\] _02467_ _04136_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_70_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09275__A2 _04593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06089__A2 _02397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08469_ _04073_ _04069_ _04074_ _04039_ _00976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_51_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10493__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10500_ _00873_ io_in[4] u_cpu.rf_ram.memory\[11\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09027__A2 _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05392__S0 _01507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10431_ _00804_ io_in[4] u_cpu.rf_ram.memory\[92\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08786__A1 u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10362_ _00009_ io_in[4] u_cpu.rf_ram_if.rdata0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05667__C _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05144__S0 _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06261__A2 _02707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10293_ _00679_ io_in[4] u_cpu.rf_ram.memory\[130\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09709__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07761__A2 _03583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05772__A1 u_cpu.cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09859__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07513__A2 _03435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05903__S _02431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05524__A1 _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10836__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09266__A2 _04593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09018__A2 _04453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07029__A1 _02642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10986__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08226__B1 _03829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10629_ _01002_ io_in[4] u_cpu.rf_ram.memory\[32\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08777__A1 _03705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07629__I _02666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05135__S0 _01522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06252__A2 _02707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10216__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08529__A1 _03935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07201__A1 _02667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07840_ _03500_ _03626_ _03629_ _00791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04988__I _01499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07752__A2 _03573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10366__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07771_ _03506_ _03583_ _03589_ _00762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_04983_ _01498_ _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_49_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09510_ _04738_ _01353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06722_ _02895_ _02988_ _02995_ _00307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07504__A2 _03435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09441_ u_cpu.rf_ram.memory\[111\]\[3\] _04691_ _04695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06653_ u_cpu.rf_ram.memory\[40\]\[0\] _02956_ _02957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05515__A1 _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05604_ u_cpu.rf_ram.memory\[0\]\[7\] u_cpu.rf_ram.memory\[1\]\[7\] u_cpu.rf_ram.memory\[2\]\[7\]
+ u_cpu.rf_ram.memory\[3\]\[7\] _01508_ _01509_ _02182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09372_ _02652_ _04651_ _04656_ _01297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09257__A2 _04583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06584_ _02464_ _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_36_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08323_ _03936_ _03950_ _03951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08465__B1 _04070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05535_ _01548_ _02113_ _01480_ _02114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_32_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05818__A2 _01467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05466_ u_cpu.rf_ram.memory\[120\]\[5\] u_cpu.rf_ram.memory\[121\]\[5\] u_cpu.rf_ram.memory\[122\]\[5\]
+ u_cpu.rf_ram.memory\[123\]\[5\] _01598_ _01556_ _02046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08254_ u_cpu.rf_ram.memory\[113\]\[2\] _03885_ _03888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09009__A2 _02870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07205_ _03098_ _03267_ _03268_ _00517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08217__B1 _03829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06491__A2 _02851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08185_ _03842_ _03843_ _00923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05397_ u_cpu.rf_ram.memory\[68\]\[4\] u_cpu.rf_ram.memory\[69\]\[4\] u_cpu.rf_ram.memory\[70\]\[4\]
+ u_cpu.rf_ram.memory\[71\]\[4\] _01507_ _01605_ _01978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08144__B _02915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07136_ u_cpu.rf_ram.memory\[53\]\[2\] _03227_ _03230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05126__S0 _01496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07067_ _03106_ _03187_ _03191_ _00456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06243__A2 _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11141__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06018_ u_arbiter.i_wb_cpu_dbus_adr\[17\] _02397_ _02523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07991__A2 _03720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10709__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07274__I _02631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07743__A2 _03573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07969_ _02965_ _03037_ _03709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09708_ _00102_ io_in[4] u_cpu.rf_ram.memory\[82\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10859__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10980_ _01349_ io_in[4] u_cpu.cpu.genblk3.csr.mcause3_0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09496__A2 _04723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09639_ _04622_ _04812_ _04813_ _01407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05506__A1 _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09248__A2 _04583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07259__A1 _02632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08456__C2 _03925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08208__B1 _03833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06482__A2 _02840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10239__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08759__A1 _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10414_ _00787_ io_in[4] u_cpu.rf_ram.memory\[91\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09420__A2 _04681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07431__A1 _03310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06234__A2 _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10345_ _00731_ io_in[4] u_cpu.rf_ram.memory\[125\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07982__A2 _03710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10389__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10276_ _00662_ io_in[4] u_cpu.rf_ram.memory\[132\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09184__A1 _04444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07734__A2 _03563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08931__A1 _03932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08931__B2 _03944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05745__A1 u_cpu.cpu.immdec.imm31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09487__A2 _02303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07498__A1 _02976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09239__A2 _04573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11014__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05320_ u_cpu.rf_ram.memory\[132\]\[3\] u_cpu.rf_ram.memory\[133\]\[3\] u_cpu.rf_ram.memory\[134\]\[3\]
+ u_cpu.rf_ram.memory\[135\]\[3\] _01634_ _01635_ _01902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_119_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05356__S0 _01496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05251_ _01493_ _01832_ _01833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06473__A2 _02840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05182_ u_cpu.rf_ram.memory\[56\]\[2\] u_cpu.rf_ram.memory\[57\]\[2\] u_cpu.rf_ram.memory\[58\]\[2\]
+ u_cpu.rf_ram.memory\[59\]\[2\] _01567_ _01568_ _01765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09411__A2 _04671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05659__S1 _01622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06225__A2 _02679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05100__C _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09990_ _00384_ io_in[4] u_cpu.rf_ram.memory\[64\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08470__I0 u_arbiter.i_wb_cpu_rdt\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07973__A2 _03710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08941_ _03986_ _03949_ _03965_ _04403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08872_ _02731_ _02825_ _04360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_57_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07725__A2 _03563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07823_ u_cpu.rf_ram.memory\[91\]\[3\] _03616_ _03620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05736__A1 _01445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05051__I3 u_cpu.rf_ram.memory\[139\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07754_ u_cpu.rf_ram.memory\[38\]\[6\] _03573_ _03580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04966_ _01495_ _01551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09478__A2 _04711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08525__I1 u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07489__A1 _03314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06705_ u_cpu.rf_ram.memory\[129\]\[7\] _02978_ _02986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07685_ _03510_ _03533_ _03541_ _00724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_04897_ u_cpu.cpu.immdec.imm24_20\[2\] _01469_ _01484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08150__A2 _02915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09424_ _04630_ _04681_ _04685_ _01320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_64_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06636_ u_cpu.rf_ram.memory\[17\]\[1\] _02945_ _02947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06161__A1 _02628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05595__S0 _01522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09355_ u_cpu.rf_ram.memory\[59\]\[5\] _04641_ _04647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06567_ _02899_ _02900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_100_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08306_ _02466_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[12\] _03934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05518_ u_cpu.rf_ram.memory\[8\]\[6\] u_cpu.rf_ram.memory\[9\]\[6\] u_cpu.rf_ram.memory\[10\]\[6\]
+ u_cpu.rf_ram.memory\[11\]\[6\] _01497_ _01525_ _02097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09286_ _04438_ _04603_ _04605_ _01262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05347__S0 _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06498_ _02689_ _02851_ _02857_ _00221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09650__A2 _04812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07661__A1 _03504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08237_ u_arbiter.i_wb_cpu_rdt\[27\] _03807_ _03829_ u_arbiter.i_wb_cpu_dbus_dat\[28\]
+ _03878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06464__A2 _02829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05449_ _01571_ _02028_ _02029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08168_ _03830_ _03831_ _00918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09402__A2 _04671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10531__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06216__A2 _02679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07119_ _03104_ _03217_ _03220_ _00479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07413__A1 _03310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08099_ u_cpu.rf_ram.memory\[116\]\[1\] _03780_ _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07964__A2 _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10130_ _00007_ io_in[4] u_cpu.rf_ram.rdata\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09166__A1 _04444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10061_ _00455_ io_in[4] u_cpu.rf_ram.memory\[57\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10681__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08913__A1 _03695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07716__A2 _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05727__A1 u_cpu.cpu.state.genblk1.misalign_trap_sync_r vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09469__A2 _02954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11037__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10963_ _01332_ io_in[4] u_cpu.rf_ram.memory\[111\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08141__A2 _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10894_ _01263_ io_in[4] u_cpu.rf_ram.memory\[108\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05586__S0 _01523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10061__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05338__S0 _01523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09641__A2 _04812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06455__A2 _02829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06207__A2 _02679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07955__A2 _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10328_ _00714_ io_in[4] u_cpu.rf_ram.memory\[127\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05966__A1 _02418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10259_ _00645_ io_in[4] u_cpu.rf_ram.memory\[134\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07707__A2 _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08904__A1 u_cpu.rf_ram.memory\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05718__A1 u_cpu.cpu.state.o_cnt_r\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06391__A1 _02669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05590__C _01466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08132__A2 _02355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10404__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07470_ u_cpu.rf_ram.memory\[136\]\[3\] _03415_ _03419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05577__S0 _01529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06421_ u_cpu.rf_ram.memory\[45\]\[6\] _02805_ _02812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06694__A2 _02978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09140_ _04434_ _04523_ _04524_ _01197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06352_ u_cpu.rf_ram.memory\[78\]\[1\] _02770_ _02772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05329__S0 _01497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09632__A2 _04802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05303_ _01602_ _01884_ _01885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10554__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09071_ u_arbiter.i_wb_cpu_rdt\[17\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\]
+ _04485_ _04487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06283_ u_cpu.cpu.immdec.imm11_7\[2\] _02728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07643__A1 _03504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08840__B1 _04329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08022_ _02667_ _03730_ _03738_ _00865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05234_ u_cpu.rf_ram.memory\[128\]\[2\] u_cpu.rf_ram.memory\[129\]\[2\] u_cpu.rf_ram.memory\[130\]\[2\]
+ u_cpu.rf_ram.memory\[131\]\[2\] _01641_ _01642_ _01817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09396__A1 _04638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08199__A2 _03822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05165_ _01528_ _01747_ _01534_ _01748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__04950__B _01534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08422__B _04039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07946__A2 _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09973_ _00367_ io_in[4] u_cpu.rf_ram.memory\[66\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05096_ u_cpu.rf_ram.memory\[52\]\[1\] u_cpu.rf_ram.memory\[53\]\[1\] u_cpu.rf_ram.memory\[54\]\[1\]
+ u_cpu.rf_ram.memory\[55\]\[1\] _01572_ _01573_ _01680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__05957__A1 _02389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09148__A1 _04444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08924_ u_cpu.rf_ram.memory\[93\]\[7\] _04381_ _04389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08746__I1 u_arbiter.i_wb_cpu_dbus_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08855_ _04350_ _04351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08371__A2 _03956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07806_ _03609_ _02927_ _03610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_57_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08786_ u_arbiter.i_wb_cpu_ibus_adr\[1\] _04309_ _04311_ u_cpu.cpu.ctrl.o_ibus_adr\[2\]
+ _04313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05998_ u_cpu.cpu.ctrl.o_ibus_adr\[12\] _02499_ u_cpu.cpu.ctrl.o_ibus_adr\[13\] _02507_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_26_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07737_ _03508_ _03563_ _03570_ _00747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04949_ _01519_ _01534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08123__A2 _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10084__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07668_ _02766_ _02965_ _03532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05568__S0 _01507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09407_ u_cpu.rf_ram.memory\[110\]\[4\] _04671_ _04676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06619_ _02885_ _02935_ _02937_ _00262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07882__A1 _03504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06685__A2 _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07599_ _02652_ _03485_ _03490_ _00689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09338_ u_cpu.rf_ram.memory\[84\]\[6\] _04624_ _04637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09623__A2 _04802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06437__A2 _02816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07634__A1 u_cpu.rf_ram.memory\[128\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09269_ u_cpu.rf_ram.memory\[83\]\[2\] _04593_ _04596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04999__A2 _01521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07937__A2 _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11162_ io_oeb[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_122_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05948__A1 _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10113_ _00507_ io_in[4] u_cpu.rf_ram.memory\[9\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11093_ _00081_ io_in[0] u_arbiter.i_wb_cpu_rdt\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10044_ _00438_ io_in[4] u_cpu.rf_ram.memory\[5\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08362__A2 _03908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05691__B u_cpu.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10427__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06373__A1 _02669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10946_ _01315_ io_in[4] u_cpu.rf_ram.memory\[110\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06125__A1 u_cpu.cpu.decode.op26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05911__S _02431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10577__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06676__A2 _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10877_ _01246_ io_in[4] u_cpu.rf_ram.memory\[107\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05710__I u_cpu.cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09614__A2 _04792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07625__A1 _03506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06428__A2 _02816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08822__B1 _04329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05100__A2 _01679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09378__A1 _02667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07928__A2 _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08050__A1 _03699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06600__A2 _02397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06970_ u_cpu.rf_ram.memory\[61\]\[0\] _03137_ _03138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05921_ _02447_ _00052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08640_ _02305_ _02320_ _04227_ _04228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_66_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05852_ _02355_ _02407_ _02408_ _02409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__04996__I _01485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05167__A2 _01749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08571_ _04143_ _04165_ _04166_ _04019_ _00986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_82_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05783_ _02353_ _02354_ _02357_ _00798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_54_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08105__A2 _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09302__A1 _04434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07522_ u_cpu.rf_ram.memory\[133\]\[2\] _03445_ _03448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05106__B _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06116__A1 _01460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07864__A1 _02286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07453_ _03314_ _03405_ _03409_ _00624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06667__A2 _02956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06404_ u_cpu.rf_ram.memory\[46\]\[7\] _02794_ _02802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07384_ u_cpu.rf_ram.memory\[14\]\[5\] _03365_ _03371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09605__A2 _04792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09123_ u_cpu.rf_ram.memory\[102\]\[1\] _04513_ _04515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07616__A1 _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06419__A2 _02805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06335_ _02685_ _02756_ _02760_ _00155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09054_ u_cpu.rf_ram.memory\[28\]\[1\] _04476_ _04478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06266_ _02718_ _02719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07092__A2 _03197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08005_ _02731_ _02954_ _03729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05217_ _01617_ _01799_ _01607_ _01800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_132_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06197_ _02609_ _02673_ _02674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07919__A2 _03672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08041__A1 _02754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05148_ u_cpu.rf_ram.memory\[140\]\[1\] u_cpu.rf_ram.memory\[141\]\[1\] u_cpu.rf_ram.memory\[142\]\[1\]
+ u_cpu.rf_ram.memory\[143\]\[1\] _01641_ _01642_ _01732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_116_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08592__A2 _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05079_ _01528_ _01662_ _01663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09956_ _00350_ io_in[4] u_cpu.rf_ram.memory\[68\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08907_ _02667_ _04371_ _04379_ _01109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09887_ _00281_ io_in[4] u_cpu.rf_ram.memory\[40\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09742__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09541__A1 _04634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08344__A2 _03938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08838_ u_cpu.cpu.ctrl.o_ibus_adr\[26\] _04327_ _04329_ u_cpu.cpu.ctrl.o_ibus_adr\[27\]
+ _04340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06355__A1 _02683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05158__A2 _01740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07282__I _02641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08769_ _03697_ _04299_ _04302_ _01048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10800_ _01169_ io_in[4] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05016__B _01600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09892__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10731_ _01100_ io_in[4] u_cpu.rf_ram.memory\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06658__A2 _02956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07855__A1 u_cpu.cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10662_ _01035_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05330__A2 _01910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07607__A1 _02677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08804__B1 _04311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10593_ _00966_ io_in[4] u_cpu.rf_ram.memory\[114\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08280__A1 _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07083__A2 _03197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06830__A2 _03049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08032__A1 _02647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11145_ _00078_ io_in[0] u_scanchain_local.module_data_in\[57\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06594__A1 u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11076_ _01435_ io_in[4] u_cpu.rf_ram_if.rcnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08335__A2 _03906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10027_ _00421_ io_in[4] u_cpu.rf_ram.memory\[60\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06346__A1 _02728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06897__A2 _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07846__A1 _03506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06649__A2 _02945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10929_ _01298_ io_in[4] u_cpu.rf_ram.memory\[10\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05321__A2 _01902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09599__A1 _04638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06120_ _01460_ _02605_ _02392_ u_cpu.cpu.o_wen0 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_117_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08271__A1 _02465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07074__A2 _03187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05596__B _01481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06051_ u_arbiter.i_wb_cpu_dbus_adr\[23\] _02397_ _02550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06821__A2 _03049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05180__S1 _01563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05002_ u_cpu.rf_ram.memory\[96\]\[0\] u_cpu.rf_ram.memory\[97\]\[0\] u_cpu.rf_ram.memory\[98\]\[0\]
+ u_cpu.rf_ram.memory\[99\]\[0\] _01567_ _01568_ _01587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__05880__I0 u_arbiter.i_wb_cpu_rdt\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08023__A1 _02731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09071__I0 u_arbiter.i_wb_cpu_rdt\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09810_ _00204_ io_in[4] u_cpu.rf_ram.memory\[51\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09765__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08574__A2 _04165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09741_ _00135_ io_in[4] u_cpu.rf_ram.memory\[20\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06953_ _03098_ _03127_ _03128_ _00405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10742__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05904_ _02438_ _00043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09672_ _02677_ _02743_ _04831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06884_ u_cpu.rf_ram.memory\[65\]\[6\] _03079_ _03086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06337__A1 _02687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08623_ _03923_ _04178_ _03910_ _04212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_36_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05835_ io_in[1] _02395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06888__A2 _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08554_ _03925_ _03998_ _04150_ _03908_ _04151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_70_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10892__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05766_ _02333_ _02334_ _02340_ _02341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_54_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05560__A2 _02134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07505_ _03312_ _03435_ _03438_ _00647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08485_ _03922_ _03908_ _03909_ _04088_ _04031_ _04089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_51_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05697_ u_cpu.rf_ram.rdata\[0\] _02273_ _02274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08147__B _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07436_ u_cpu.rf_ram.memory\[137\]\[4\] _03395_ _03400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05312__A2 _01893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10122__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07367_ _03318_ _03355_ _03361_ _00586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09106_ _04438_ _04503_ _04505_ _01182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06318_ _02652_ _02745_ _02750_ _00148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07065__A2 _03187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07298_ u_cpu.rf_ram.memory\[72\]\[7\] _03308_ _03323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09037_ u_cpu.rf_ram.memory\[96\]\[4\] _04463_ _04468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06249_ u_cpu.rf_ram.memory\[18\]\[1\] _02707_ _02709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06812__A2 _03039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10272__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05171__S1 _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08014__A1 _02647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08565__A2 _02259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05379__A2 _01959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09939_ _00333_ io_in[4] u_cpu.rf_ram.memory\[75\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06879__A2 _03079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05551__A2 _02125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07828__A1 _03506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10714_ _01084_ io_in[4] u_cpu.cpu.ctrl.o_ibus_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05303__A2 _01884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06500__A1 _02691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10645_ _01018_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10615__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08253__A1 _03695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07056__A2 _03177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10576_ _00949_ io_in[4] u_cpu.rf_ram.memory\[113\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09788__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06803__A2 _03039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05162__S1 _01525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08005__A1 _02731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10765__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08556__A2 _04000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11128_ _00060_ io_in[0] u_scanchain_local.module_data_in\[40\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08308__A2 _03935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11059_ _01427_ io_in[4] u_cpu.rf_ram.memory\[23\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05790__A2 _02265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05620_ u_cpu.rf_ram.memory\[60\]\[7\] u_cpu.rf_ram.memory\[61\]\[7\] u_cpu.rf_ram.memory\[62\]\[7\]
+ u_cpu.rf_ram.memory\[63\]\[7\] _01496_ _01594_ _02198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_24_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05542__A2 _02092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10145__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05551_ _02123_ _02125_ _02127_ _02129_ _01560_ _02130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_60_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08270_ _02465_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[2\] _03898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05482_ _02055_ _02057_ _02059_ _02061_ _01486_ _02062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__08492__A1 _04000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07295__A2 _03308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07221_ _03276_ _03277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10295__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08244__A1 u_arbiter.i_wb_cpu_rdt\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07152_ u_cpu.rf_ram.memory\[52\]\[1\] _03237_ _03239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07047__A2 _03177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06103_ _02590_ _02592_ _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07083_ _03104_ _03197_ _03200_ _00463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05153__S1 _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06034_ u_cpu.cpu.ctrl.o_ibus_adr\[20\] _02531_ _02536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_133_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06007__B1 _02398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07985_ u_cpu.rf_ram.memory\[118\]\[7\] _03710_ _03718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09724_ _00118_ io_in[4] u_cpu.rf_ram.memory\[81\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06936_ u_cpu.rf_ram.memory\[63\]\[1\] _03117_ _03119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09655_ _04821_ _04822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06867_ _02895_ _03069_ _03076_ _00371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08606_ _03912_ _04185_ _04196_ _03896_ _04197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_05818_ u_cpu.rf_ram_if.rdata0\[3\] _01467_ _02383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09586_ u_cpu.rf_ram.memory\[24\]\[1\] _04782_ _04784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06730__A1 _02885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06798_ _02731_ _03037_ _03038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05533__A2 _02111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04967__S1 _01524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08537_ _04134_ _04135_ _00983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11070__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05749_ _02322_ _02323_ _02319_ _02324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_70_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10638__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08483__A1 _03922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08468_ u_cpu.cpu.immdec.imm24_20\[3\] _04068_ _03896_ _04074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07286__A2 _03308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08483__B2 _03940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05297__A1 _01490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07419_ _03316_ _03385_ _03390_ _00609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08399_ _04009_ _04010_ _04018_ _04019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09930__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05392__S1 _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08605__B _03912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10430_ _00803_ io_in[4] u_cpu.rf_ram.memory\[92\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07038__A2 _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10788__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08786__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10361_ _00008_ io_in[4] u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05144__S1 _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10292_ _00678_ io_in[4] u_cpu.rf_ram.memory\[130\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10018__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07210__A2 _03267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10168__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08171__B1 _03833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06721__A1 u_cpu.rf_ram.memory\[139\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05080__S0 _01530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07277__A2 _03308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07029__A2 _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08226__A1 u_arbiter.i_wb_cpu_rdt\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10628_ _01001_ io_in[4] u_cpu.rf_ram.memory\[32\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08226__B2 u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08777__A2 _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10559_ _00932_ io_in[4] u_arbiter.i_wb_cpu_dbus_dat\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05135__S1 _01622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06788__A1 _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05460__A1 _01512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08529__A2 _03974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07201__A2 _03257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07770_ u_cpu.rf_ram.memory\[37\]\[5\] _03583_ _03589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04982_ _01494_ _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09803__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06721_ u_cpu.rf_ram.memory\[139\]\[6\] _02988_ _02995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11093__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09440_ _04628_ _04691_ _04694_ _01327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06652_ _02955_ _02956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05515__A2 _02093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06712__A1 _02885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05071__S0 _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05603_ _01493_ _02180_ _02181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09371_ u_cpu.rf_ram.memory\[10\]\[4\] _04651_ _04656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06583_ _02667_ _02900_ _02908_ _00255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09953__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08322_ _03939_ _03949_ _03950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05534_ u_cpu.rf_ram.memory\[56\]\[6\] u_cpu.rf_ram.memory\[57\]\[6\] u_cpu.rf_ram.memory\[58\]\[6\]
+ u_cpu.rf_ram.memory\[59\]\[6\] _01567_ _01568_ _02113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_33_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07268__A2 _03297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08465__B2 u_cpu.cpu.immdec.imm24_20\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08253_ _03695_ _03885_ _03887_ _00947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05465_ _01543_ _02044_ _02045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10930__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07204_ u_cpu.rf_ram.memory\[142\]\[0\] _03267_ _03268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08217__A1 u_arbiter.i_wb_cpu_rdt\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08184_ u_arbiter.i_wb_cpu_rdt\[9\] _03822_ _03833_ u_arbiter.i_wb_cpu_dbus_dat\[10\]
+ _03843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08217__B2 u_arbiter.i_wb_cpu_dbus_dat\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05396_ _01621_ _01976_ _01977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08768__A2 _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07135_ _03102_ _03227_ _03229_ _00486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06779__A1 _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05126__S1 _01594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07066_ u_cpu.rf_ram.memory\[57\]\[3\] _03187_ _03191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07440__A2 _03395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05451__A1 _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06017_ u_cpu.cpu.ctrl.o_ibus_adr\[17\] _02519_ _02521_ _02461_ _02522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__05784__B _01444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09193__A2 _04553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10310__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05203__A1 _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07968_ _03707_ _03693_ _03708_ _00841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_47_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06919_ _03106_ _03100_ _03107_ _00392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09707_ _00101_ io_in[4] u_cpu.rf_ram.memory\[82\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05008__C _01560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07899_ u_cpu.rf_ram.memory\[35\]\[4\] _03662_ _03667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09638_ u_cpu.rf_ram.memory\[100\]\[0\] _04812_ _04813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10460__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09569_ _04626_ _04772_ _04774_ _01376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08456__A1 _03974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07259__A2 _03297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08456__B2 _04050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08208__A1 u_arbiter.i_wb_cpu_rdt\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05678__C _01466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10413_ _00786_ io_in[4] u_cpu.rf_ram.memory\[91\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05690__A1 u_arbiter.i_wb_cpu_dbus_we vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10344_ _00730_ io_in[4] u_cpu.rf_ram.memory\[125\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07431__A2 _03395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05442__A1 _01463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10275_ _00661_ io_in[4] u_cpu.rf_ram.memory\[132\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05993__A2 _02499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09826__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09184__A2 _04543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07195__A1 _02652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08931__A2 _03975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10803__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09976__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07498__A2 _03037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10953__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08447__A1 _04024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08998__A2 _04436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05356__S1 _01594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05250_ u_cpu.rf_ram.memory\[4\]\[3\] u_cpu.rf_ram.memory\[5\]\[3\] u_cpu.rf_ram.memory\[6\]\[3\]
+ u_cpu.rf_ram.memory\[7\]\[3\] _01523_ _01525_ _01832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_80_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07670__A2 _03533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05181_ _01464_ _01763_ _01764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07422__A2 _03385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10333__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08470__I1 u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05433__A1 _01513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08940_ _04399_ _04402_ _01119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09175__A2 _04543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08871_ _03707_ _04351_ _04359_ _01093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07822_ _03500_ _03616_ _03619_ _00783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08922__A2 _04381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10483__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05736__A2 _02265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05292__S0 _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07753_ _03506_ _03573_ _03579_ _00754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_04965_ _01548_ _01549_ _01518_ _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_49_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06704_ _02895_ _02978_ _02985_ _00299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_93_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07684_ u_cpu.rf_ram.memory\[126\]\[7\] _03533_ _03541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07489__A2 _03425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08686__A1 _03707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04896_ u_cpu.cpu.immdec.imm19_12_20\[6\] _01438_ _01483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09423_ u_cpu.rf_ram.memory\[86\]\[3\] _04681_ _04685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05044__S0 _01529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06635_ _02881_ _02945_ _02946_ _00269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06161__A2 _02642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05595__S1 _01622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09354_ _04632_ _04641_ _04646_ _01289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08438__A1 _03705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06566_ _02717_ _02731_ _02899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08305_ _03926_ _03932_ _03933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_33_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08989__A2 _04436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05517_ _01528_ _02095_ _01534_ _02096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09285_ u_cpu.rf_ram.memory\[108\]\[1\] _04603_ _04605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06497_ u_cpu.rf_ram.memory\[43\]\[5\] _02851_ _02857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05347__S1 _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08236_ u_arbiter.i_wb_cpu_dbus_dat\[27\] _03808_ _03877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05448_ u_cpu.rf_ram.memory\[52\]\[5\] u_cpu.rf_ram.memory\[53\]\[5\] u_cpu.rf_ram.memory\[54\]\[5\]
+ u_cpu.rf_ram.memory\[55\]\[5\] _01572_ _01573_ _02028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07661__A2 _03523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08167_ u_arbiter.i_wb_cpu_rdt\[4\] _03822_ _03808_ u_arbiter.i_wb_cpu_dbus_dat\[4\]
+ _03831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05379_ _01597_ _01959_ _01600_ _01960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09849__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07118_ u_cpu.rf_ram.memory\[54\]\[2\] _03217_ _03220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08098_ _03691_ _03780_ _03781_ _00898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07413__A2 _03385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05424__A1 _01506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07049_ _03106_ _03177_ _03181_ _00448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10826__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05975__A2 _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07285__I _02646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09166__A2 _04533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10060_ _00454_ io_in[4] u_cpu.rf_ram.memory\[57\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07177__A1 _02652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09999__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08913__A2 _04381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05283__S0 _01529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10976__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10962_ _01331_ io_in[4] u_cpu.rf_ram.memory\[111\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10893_ _01262_ io_in[4] u_cpu.rf_ram.memory\[108\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10206__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05586__S1 _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05338__S1 _01525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07101__A1 _03104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07652__A2 _03523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10356__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05909__S _02431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08601__A1 _03928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07404__A2 _03375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05415__A1 _01986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10327_ _00713_ io_in[4] u_cpu.rf_ram.memory\[127\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09157__A2 _04533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10258_ _00644_ io_in[4] u_cpu.rf_ram.memory\[135\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08904__A2 _04371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10189_ _00575_ io_in[4] u_cpu.rf_ram.memory\[70\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05718__A2 _02290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05274__S0 _01576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06391__A2 _02794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08668__A1 _03707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05026__S0 _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05577__S1 _01500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06420_ _02689_ _02805_ _02811_ _00189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11131__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07891__A2 _03662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06351_ _02669_ _02770_ _02771_ _00160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05329__S1 _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05302_ u_cpu.rf_ram.memory\[80\]\[3\] u_cpu.rf_ram.memory\[81\]\[3\] u_cpu.rf_ram.memory\[82\]\[3\]
+ u_cpu.rf_ram.memory\[83\]\[3\] _01544_ _01594_ _01884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09070_ _04486_ _01165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06282_ _02693_ _02719_ _02727_ _00135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08690__S _04257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07643__A2 _03513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08021_ u_cpu.rf_ram.memory\[8\]\[7\] _03730_ _03738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05233_ _01638_ _01815_ _01534_ _01816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05111__C _01560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10849__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09396__A2 _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05164_ u_cpu.rf_ram.memory\[0\]\[2\] u_cpu.rf_ram.memory\[1\]\[2\] u_cpu.rf_ram.memory\[2\]\[2\]
+ u_cpu.rf_ram.memory\[3\]\[2\] _01530_ _01532_ _01747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_116_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09972_ _00366_ io_in[4] u_cpu.rf_ram.memory\[66\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05095_ _01566_ _01678_ _01480_ _01679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09148__A2 _04523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08923_ _03705_ _04381_ _04388_ _01116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10999__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07159__A1 _03108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08356__B1 _03912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08854_ _02803_ _04349_ _04350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05265__S0 _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07805_ u_cpu.rf_ram_if.rgnt _03609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_85_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08785_ _04312_ _01054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_05997_ _02389_ _02505_ _02506_ _00071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_57_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06382__A2 _02784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10229__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07736_ u_cpu.rf_ram.memory\[123\]\[6\] _03563_ _03570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04948_ u_cpu.rf_ram.memory\[0\]\[0\] u_cpu.rf_ram.memory\[1\]\[0\] u_cpu.rf_ram.memory\[2\]\[0\]
+ u_cpu.rf_ram.memory\[3\]\[0\] _01530_ _01532_ _01533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_72_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05590__B1 _02166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09320__A2 _04624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07667_ _03510_ _03523_ _03531_ _00716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04879_ u_cpu.rf_ram_if.rtrig0 _01452_ _01466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__05568__S1 _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07331__A1 _03318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09406_ _04630_ _04671_ _04675_ _01312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06618_ u_cpu.rf_ram.memory\[16\]\[1\] _02935_ _02937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07882__A2 _03652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07598_ u_cpu.rf_ram.memory\[12\]\[4\] _03485_ _03490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_90_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10379__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06549_ u_cpu.rf_ram.memory\[50\]\[2\] _02883_ _02888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09337_ _02661_ _04636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09268_ _04438_ _04593_ _04595_ _01254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07634__A2 _03513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05645__A1 _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08219_ u_arbiter.i_wb_cpu_dbus_dat\[21\] _03808_ _03866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09199_ u_cpu.rf_ram.memory\[79\]\[3\] _04553_ _04557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__04999__A3 _01542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09387__A2 _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11161_ io_oeb[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_1_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09139__A2 _04523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10112_ _00506_ io_in[4] u_cpu.rf_ram.memory\[9\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06070__A1 _02562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11092_ _00070_ io_in[0] u_arbiter.i_wb_cpu_rdt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11004__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10043_ _00437_ io_in[4] u_cpu.rf_ram.memory\[5\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05256__S0 _01530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06373__A2 _02784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07570__A1 _02619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11154__CLK io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09311__A2 _04613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10945_ _01314_ io_in[4] u_cpu.rf_ram.memory\[110\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06125__A2 u_cpu.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10876_ _01245_ io_in[4] u_cpu.rf_ram.memory\[107\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07873__A2 _03652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07625__A2 _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05636__A1 _01512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09378__A2 _04651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07389__A1 _02667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08050__A2 _03750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05920_ u_arbiter.i_wb_cpu_rdt\[30\] u_arbiter.i_wb_cpu_dbus_dat\[27\] _02431_ _02447_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08889__A1 _02667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05247__S0 _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09550__A2 _04762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05851_ _01441_ _02402_ _02408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06364__A2 _02770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07561__A1 _03314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08570_ u_cpu.cpu.immdec.imm19_12_20\[1\] _03897_ _04165_ _04166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05782_ _02354_ _02356_ _02357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07521_ _03310_ _03445_ _03447_ _00654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09302__A2 _04613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10521__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07313__A1 _03318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07452_ u_cpu.rf_ram.memory\[49\]\[3\] _03405_ _03409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06403_ _02691_ _02794_ _02801_ _00182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07383_ _02652_ _03365_ _03370_ _00593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09122_ _04434_ _04513_ _04514_ _01189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10671__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06334_ u_cpu.rf_ram.memory\[80\]\[3\] _02756_ _02760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07616__A2 _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05627__A1 _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09053_ _04434_ _04476_ _04477_ _01157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06265_ _02677_ _02717_ _02718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08004_ _03707_ _03720_ _03728_ _00857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05216_ u_cpu.rf_ram.memory\[84\]\[2\] u_cpu.rf_ram.memory\[85\]\[2\] u_cpu.rf_ram.memory\[86\]\[2\]
+ u_cpu.rf_ram.memory\[87\]\[2\] _01507_ _01605_ _01799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09369__A2 _04651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06196_ _01460_ _02610_ _02612_ _02673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__11027__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05147_ _01465_ _01730_ _01731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08041__A2 _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09955_ _00349_ io_in[4] u_cpu.rf_ram.memory\[68\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05078_ u_cpu.rf_ram.memory\[8\]\[1\] u_cpu.rf_ram.memory\[9\]\[1\] u_cpu.rf_ram.memory\[10\]\[1\]
+ u_cpu.rf_ram.memory\[11\]\[1\] _01523_ _01525_ _01662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_106_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08906_ u_cpu.rf_ram.memory\[2\]\[7\] _04371_ _04379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10051__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09886_ _00280_ io_in[4] u_cpu.rf_ram.memory\[40\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09541__A2 _04752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08837_ _04339_ _01079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_44_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06355__A2 _02770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07552__A1 _02825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08768_ u_cpu.rf_ram.memory\[30\]\[2\] _04299_ _04302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07719_ _03508_ _03553_ _03560_ _00739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08699_ _04262_ _01018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_81_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10730_ _01099_ io_in[4] u_cpu.rf_ram.memory\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07855__A2 _01442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08327__C _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05410__S0 _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09057__A1 _04440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10661_ _01034_ io_in[4] u_arbiter.i_wb_cpu_dbus_adr\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07607__A2 _03037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10592_ _00965_ io_in[4] u_cpu.rf_ram.memory\[114\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05618__A1 _01463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08280__A2 u_arbiter.i_wb_cpu_rdt\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08032__A2 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11144_ _00077_ io_in[0] u_scanchain_local.module_data_in\[56\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07791__A1 _03508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11075_ u_cpu.rf_ram_if.rtrig0 io_in[4] u_cpu.rf_ram_if.rtrig1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08569__I _04164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10026_ _00420_ io_in[4] u_cpu.rf_ram.memory\[61\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09532__A2 _04752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10544__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07543__A1 _03314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06346__A2 _02608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05207__B _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05922__S _02431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09296__A1 _04448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08099__A2 _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10694__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07846__A2 _03626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10928_ _01297_ io_in[4] u_cpu.rf_ram.memory\[10\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05401__S0 _01529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09048__A1 _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10859_ _01228_ io_in[4] u_cpu.rf_ram.memory\[79\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09599__A2 _04782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05609__A1 _01464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08271__A2 _02414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06282__A1 _02693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06050_ _02461_ _02548_ _02549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05001_ _01571_ _01585_ _01586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05880__I1 u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10074__CLK io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09220__A1 _04444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08023__A2 _02849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05468__S0 _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06585__A2 _02461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09740_ _00134_ io_in[4] u_cpu.rf_ram.memory\[20\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06952_ u_cpu.rf_ram.memory\[62\]\[0\] _03127_ _03128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
.ends

