magic
tech gf180mcuC
magscale 1 5
timestamp 1670234014
<< obsm1 >>
rect 672 1538 99288 58438
<< obsm2 >>
rect 910 233 99778 58427
<< metal3 >>
rect 99800 57792 100000 57848
rect 99800 53816 100000 53872
rect 99800 49840 100000 49896
rect 99800 45864 100000 45920
rect 99800 41888 100000 41944
rect 99800 37912 100000 37968
rect 99800 33936 100000 33992
rect 99800 29960 100000 30016
rect 99800 25984 100000 26040
rect 99800 22008 100000 22064
rect 99800 18032 100000 18088
rect 99800 14056 100000 14112
rect 99800 10080 100000 10136
rect 99800 6104 100000 6160
rect 99800 2128 100000 2184
<< obsm3 >>
rect 905 57878 99800 58422
rect 905 57762 99770 57878
rect 905 53902 99800 57762
rect 905 53786 99770 53902
rect 905 49926 99800 53786
rect 905 49810 99770 49926
rect 905 45950 99800 49810
rect 905 45834 99770 45950
rect 905 41974 99800 45834
rect 905 41858 99770 41974
rect 905 37998 99800 41858
rect 905 37882 99770 37998
rect 905 34022 99800 37882
rect 905 33906 99770 34022
rect 905 30046 99800 33906
rect 905 29930 99770 30046
rect 905 26070 99800 29930
rect 905 25954 99770 26070
rect 905 22094 99800 25954
rect 905 21978 99770 22094
rect 905 18118 99800 21978
rect 905 18002 99770 18118
rect 905 14142 99800 18002
rect 905 14026 99770 14142
rect 905 10166 99800 14026
rect 905 10050 99770 10166
rect 905 6190 99800 10050
rect 905 6074 99770 6190
rect 905 2214 99800 6074
rect 905 2098 99770 2214
rect 905 238 99800 2098
<< metal4 >>
rect 2224 1538 2384 58438
rect 9904 1538 10064 58438
rect 17584 1538 17744 58438
rect 25264 1538 25424 58438
rect 32944 1538 33104 58438
rect 40624 1538 40784 58438
rect 48304 1538 48464 58438
rect 55984 1538 56144 58438
rect 63664 1538 63824 58438
rect 71344 1538 71504 58438
rect 79024 1538 79184 58438
rect 86704 1538 86864 58438
rect 94384 1538 94544 58438
<< obsm4 >>
rect 4214 1508 9874 56607
rect 10094 1508 17554 56607
rect 17774 1508 25234 56607
rect 25454 1508 32914 56607
rect 33134 1508 40594 56607
rect 40814 1508 48274 56607
rect 48494 1508 55954 56607
rect 56174 1508 63634 56607
rect 63854 1508 71314 56607
rect 71534 1508 78994 56607
rect 79214 1508 86674 56607
rect 86894 1508 94354 56607
rect 94574 1508 99050 56607
rect 4214 289 99050 1508
<< labels >>
rlabel metal3 s 99800 2128 100000 2184 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 99800 6104 100000 6160 6 io_in[1]
port 2 nsew signal input
rlabel metal3 s 99800 10080 100000 10136 6 io_in[2]
port 3 nsew signal input
rlabel metal3 s 99800 14056 100000 14112 6 io_in[3]
port 4 nsew signal input
rlabel metal3 s 99800 18032 100000 18088 6 io_in[4]
port 5 nsew signal input
rlabel metal3 s 99800 41888 100000 41944 6 io_oeb[0]
port 6 nsew signal output
rlabel metal3 s 99800 45864 100000 45920 6 io_oeb[1]
port 7 nsew signal output
rlabel metal3 s 99800 49840 100000 49896 6 io_oeb[2]
port 8 nsew signal output
rlabel metal3 s 99800 53816 100000 53872 6 io_oeb[3]
port 9 nsew signal output
rlabel metal3 s 99800 57792 100000 57848 6 io_oeb[4]
port 10 nsew signal output
rlabel metal3 s 99800 22008 100000 22064 6 io_out[0]
port 11 nsew signal output
rlabel metal3 s 99800 25984 100000 26040 6 io_out[1]
port 12 nsew signal output
rlabel metal3 s 99800 29960 100000 30016 6 io_out[2]
port 13 nsew signal output
rlabel metal3 s 99800 33936 100000 33992 6 io_out[3]
port 14 nsew signal output
rlabel metal3 s 99800 37912 100000 37968 6 io_out[4]
port 15 nsew signal output
rlabel metal4 s 2224 1538 2384 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 58438 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 58438 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 58438 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 58438 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 58438 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 58438 6 vss
port 17 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 100000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 17924888
string GDS_FILE /home/runner/work/gf180-mpw0-serv/gf180-mpw0-serv/openlane/serv_1/runs/22_12_05_09_48/results/signoff/serv_1.magic.gds
string GDS_START 350324
<< end >>

