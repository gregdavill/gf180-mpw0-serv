VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO serv_1
  CLASS BLOCK ;
  FOREIGN serv_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1000.000 BY 600.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 998.000 21.280 1000.000 21.840 ;
    END
  END io_in[0]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 998.000 61.040 1000.000 61.600 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 998.000 100.800 1000.000 101.360 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 998.000 140.560 1000.000 141.120 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 998.000 180.320 1000.000 180.880 ;
    END
  END io_in[4]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 998.000 418.880 1000.000 419.440 ;
    END
  END io_oeb[0]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 998.000 458.640 1000.000 459.200 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 998.000 498.400 1000.000 498.960 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 998.000 538.160 1000.000 538.720 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 998.000 577.920 1000.000 578.480 ;
    END
  END io_oeb[4]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 998.000 220.080 1000.000 220.640 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 998.000 259.840 1000.000 260.400 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 998.000 299.600 1000.000 300.160 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 998.000 339.360 1000.000 339.920 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 998.000 379.120 1000.000 379.680 ;
    END
  END io_out[4]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 584.380 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 584.380 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 992.880 584.380 ;
      LAYER Metal2 ;
        RECT 9.100 2.330 997.780 584.270 ;
      LAYER Metal3 ;
        RECT 9.050 578.780 998.000 584.220 ;
        RECT 9.050 577.620 997.700 578.780 ;
        RECT 9.050 539.020 998.000 577.620 ;
        RECT 9.050 537.860 997.700 539.020 ;
        RECT 9.050 499.260 998.000 537.860 ;
        RECT 9.050 498.100 997.700 499.260 ;
        RECT 9.050 459.500 998.000 498.100 ;
        RECT 9.050 458.340 997.700 459.500 ;
        RECT 9.050 419.740 998.000 458.340 ;
        RECT 9.050 418.580 997.700 419.740 ;
        RECT 9.050 379.980 998.000 418.580 ;
        RECT 9.050 378.820 997.700 379.980 ;
        RECT 9.050 340.220 998.000 378.820 ;
        RECT 9.050 339.060 997.700 340.220 ;
        RECT 9.050 300.460 998.000 339.060 ;
        RECT 9.050 299.300 997.700 300.460 ;
        RECT 9.050 260.700 998.000 299.300 ;
        RECT 9.050 259.540 997.700 260.700 ;
        RECT 9.050 220.940 998.000 259.540 ;
        RECT 9.050 219.780 997.700 220.940 ;
        RECT 9.050 181.180 998.000 219.780 ;
        RECT 9.050 180.020 997.700 181.180 ;
        RECT 9.050 141.420 998.000 180.020 ;
        RECT 9.050 140.260 997.700 141.420 ;
        RECT 9.050 101.660 998.000 140.260 ;
        RECT 9.050 100.500 997.700 101.660 ;
        RECT 9.050 61.900 998.000 100.500 ;
        RECT 9.050 60.740 997.700 61.900 ;
        RECT 9.050 22.140 998.000 60.740 ;
        RECT 9.050 20.980 997.700 22.140 ;
        RECT 9.050 2.380 998.000 20.980 ;
      LAYER Metal4 ;
        RECT 42.140 15.080 98.740 566.070 ;
        RECT 100.940 15.080 175.540 566.070 ;
        RECT 177.740 15.080 252.340 566.070 ;
        RECT 254.540 15.080 329.140 566.070 ;
        RECT 331.340 15.080 405.940 566.070 ;
        RECT 408.140 15.080 482.740 566.070 ;
        RECT 484.940 15.080 559.540 566.070 ;
        RECT 561.740 15.080 636.340 566.070 ;
        RECT 638.540 15.080 713.140 566.070 ;
        RECT 715.340 15.080 789.940 566.070 ;
        RECT 792.140 15.080 866.740 566.070 ;
        RECT 868.940 15.080 943.540 566.070 ;
        RECT 945.740 15.080 990.500 566.070 ;
        RECT 42.140 2.890 990.500 15.080 ;
  END
END serv_1
END LIBRARY

