VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tiny_user_project
  CLASS BLOCK ;
  FOREIGN tiny_user_project ;
  ORIGIN 0.000 0.000 ;
  SIZE 780.000 BY 1080.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 641.760 4.000 642.320 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 651.840 4.000 652.400 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 319.200 4.000 319.760 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 561.120 4.000 561.680 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 383.040 4.000 383.600 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 329.280 4.000 329.840 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 339.360 1076.000 339.920 1079.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 336.000 779.000 336.560 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 1028.160 779.000 1028.720 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 473.760 1076.000 474.320 1079.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 131.040 779.000 131.600 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1044.960 4.000 1045.520 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 591.360 1076.000 591.920 1079.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 651.840 1.000 652.400 4.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 776.160 1076.000 776.720 1079.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 954.240 779.000 954.800 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 769.440 1.000 770.000 4.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 1.000 124.880 4.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 776.160 4.000 776.720 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 635.040 4.000 635.600 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 722.400 4.000 722.960 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 581.280 4.000 581.840 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 1071.840 779.000 1072.400 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 608.160 1.000 608.720 4.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 393.120 4.000 393.680 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 6.720 779.000 7.280 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 97.440 4.000 98.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 829.920 4.000 830.480 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 678.720 1076.000 679.280 1079.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 974.400 779.000 974.960 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 856.800 779.000 857.360 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 1061.760 779.000 1062.320 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 571.200 779.000 571.760 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 178.080 4.000 178.640 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 329.280 779.000 329.840 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 608.160 1076.000 608.720 1079.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 426.720 4.000 427.280 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 480.480 4.000 481.040 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 803.040 779.000 803.600 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 749.280 779.000 749.840 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 964.320 4.000 964.880 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 571.200 1.000 571.760 4.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 238.560 4.000 239.120 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 70.560 779.000 71.120 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 436.800 1076.000 437.360 1079.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 265.440 1.000 266.000 4.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 87.360 1.000 87.920 4.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 974.400 4.000 974.960 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 178.080 1076.000 178.640 1079.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 97.440 1076.000 98.000 1079.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 383.040 1076.000 383.600 1079.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 16.800 779.000 17.360 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 389.760 779.000 390.320 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 752.640 1076.000 753.200 1079.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 265.440 4.000 266.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 131.040 4.000 131.600 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 850.080 4.000 850.640 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 776.160 1.000 776.720 4.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 947.520 4.000 948.080 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 624.960 779.000 625.520 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 507.360 779.000 507.920 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 97.440 779.000 98.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 285.600 4.000 286.160 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 661.920 1076.000 662.480 1079.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 302.400 779.000 302.960 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 759.360 4.000 759.920 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 991.200 779.000 991.760 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 366.240 1076.000 366.800 1079.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 524.160 779.000 524.720 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 695.520 4.000 696.080 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 124.320 4.000 124.880 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 527.520 1076.000 528.080 1079.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 732.480 4.000 733.040 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 295.680 1076.000 296.240 1079.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 463.680 4.000 464.240 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 1055.040 779.000 1055.600 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1076.000 0.560 1079.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 134.400 1076.000 134.960 1079.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 598.080 1.000 598.640 4.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 759.360 1076.000 759.920 1079.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 927.360 4.000 927.920 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 688.800 4.000 689.360 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 372.960 1.000 373.520 4.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 927.360 779.000 927.920 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 104.160 1.000 104.720 4.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 87.360 779.000 87.920 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 53.760 1076.000 54.320 1079.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 60.480 1.000 61.040 4.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 238.560 779.000 239.120 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 614.880 4.000 615.440 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 356.160 779.000 356.720 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 346.080 4.000 346.640 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 33.600 779.000 34.160 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 174.720 779.000 175.280 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 393.120 1.000 393.680 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 312.480 1.000 313.040 4.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 500.640 1076.000 501.200 1079.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 635.040 1.000 635.600 4.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 480.480 779.000 481.040 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 698.880 1076.000 699.440 1079.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 329.280 1.000 329.840 4.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 430.080 1076.000 430.640 1079.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 339.360 4.000 339.920 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 614.880 1.000 615.440 4.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 554.400 1.000 554.960 4.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 221.760 1.000 222.320 4.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 43.680 4.000 44.240 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 275.520 1076.000 276.080 1079.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 426.720 1.000 427.280 4.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 241.920 1076.000 242.480 1079.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 168.000 4.000 168.560 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 527.520 4.000 528.080 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 678.720 1.000 679.280 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 238.560 1.000 239.120 4.000 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 473.760 4.000 474.320 ;
    END
  END la_data_in[0]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 1018.080 779.000 1018.640 ;
    END
  END la_data_in[10]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 561.120 779.000 561.680 ;
    END
  END la_data_in[11]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 285.600 1.000 286.160 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 221.760 1076.000 222.320 1079.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 813.120 4.000 813.680 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 819.840 779.000 820.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1018.080 4.000 1018.640 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 292.320 779.000 292.880 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 312.480 1076.000 313.040 1079.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 141.120 4.000 141.680 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 60.480 1076.000 61.040 1079.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 346.080 779.000 346.640 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 705.600 4.000 706.160 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 409.920 4.000 410.480 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 846.720 779.000 847.280 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 322.560 1076.000 323.120 1079.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 43.680 1076.000 44.240 1079.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 420.000 1076.000 420.560 1079.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 840.000 4.000 840.560 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 876.960 4.000 877.520 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 383.040 779.000 383.600 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 258.720 1076.000 259.280 1079.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 70.560 4.000 71.120 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 635.040 1076.000 635.600 1079.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 372.960 4.000 373.520 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 624.960 4.000 625.520 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1001.280 4.000 1001.840 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 823.200 4.000 823.760 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 661.920 1.000 662.480 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 910.560 4.000 911.120 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 420.000 1.000 420.560 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 356.160 1076.000 356.720 1079.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 658.560 779.000 659.120 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 319.200 1.000 319.760 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 446.880 1.000 447.440 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 312.480 4.000 313.040 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 725.760 1076.000 726.320 1079.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 157.920 779.000 158.480 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 302.400 1.000 302.960 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 829.920 779.000 830.480 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 581.280 1.000 581.840 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 285.600 1076.000 286.160 1079.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 204.960 1076.000 205.520 1079.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1008.000 4.000 1008.560 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 215.040 1076.000 215.600 1079.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 436.800 1.000 437.360 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 463.680 779.000 464.240 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 571.200 1076.000 571.760 1079.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 510.720 1076.000 511.280 1079.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 248.640 4.000 249.200 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 275.520 4.000 276.080 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 954.240 4.000 954.800 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 339.360 1.000 339.920 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 1001.280 779.000 1001.840 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 157.920 1.000 158.480 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 766.080 779.000 766.640 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 23.520 4.000 24.080 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 544.320 1.000 544.880 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 87.360 1076.000 87.920 1079.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 184.800 1.000 185.360 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 490.560 779.000 491.120 ;
    END
  END la_data_in[7]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 16.800 4.000 17.360 ;
    END
  END la_data_in[8]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 688.800 1076.000 689.360 1079.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 651.840 1076.000 652.400 1079.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 651.840 779.000 652.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 33.600 4.000 34.160 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 668.640 4.000 669.200 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 346.080 1.000 346.640 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 534.240 779.000 534.800 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 796.320 4.000 796.880 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 668.640 779.000 669.200 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 302.400 1076.000 302.960 1079.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 920.640 779.000 921.200 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 490.560 1.000 491.120 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 588.000 779.000 588.560 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 282.240 779.000 282.800 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 920.640 4.000 921.200 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 732.480 779.000 733.040 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 275.520 1.000 276.080 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 420.000 4.000 420.560 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 500.640 1.000 501.200 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 903.840 4.000 904.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 409.920 1076.000 410.480 1079.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 893.760 779.000 894.320 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 399.840 1.000 400.400 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 211.680 4.000 212.240 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 577.920 779.000 578.480 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 194.880 779.000 195.440 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 393.120 1076.000 393.680 1079.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 319.200 779.000 319.760 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 453.600 1.000 454.160 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 349.440 1076.000 350.000 1079.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 900.480 779.000 901.040 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 517.440 779.000 518.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 168.000 779.000 168.560 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 275.520 779.000 276.080 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 151.200 4.000 151.760 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 124.320 779.000 124.880 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 436.800 779.000 437.360 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 937.440 779.000 938.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 50.400 1.000 50.960 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 383.040 1.000 383.600 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1071.840 4.000 1072.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1061.760 4.000 1062.320 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 661.920 4.000 662.480 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 211.680 1.000 212.240 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 60.480 779.000 61.040 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 376.320 1076.000 376.880 1079.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 168.000 1076.000 168.560 1079.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 893.760 4.000 894.320 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 211.680 779.000 212.240 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 883.680 4.000 884.240 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 786.240 779.000 786.800 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 194.880 1076.000 195.440 1079.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 372.960 779.000 373.520 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 554.400 1076.000 554.960 1079.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 792.960 779.000 793.520 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 356.160 4.000 356.720 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 705.600 779.000 706.160 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 598.080 1076.000 598.640 1079.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 248.640 1.000 249.200 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 23.520 779.000 24.080 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 221.760 779.000 222.320 ;
    END
  END la_data_out[63]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 416.640 779.000 417.200 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 742.560 1076.000 743.120 1079.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 50.400 4.000 50.960 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 598.080 779.000 598.640 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 497.280 779.000 497.840 ;
    END
  END la_oenb[0]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 813.120 779.000 813.680 ;
    END
  END la_oenb[10]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 678.720 779.000 679.280 ;
    END
  END la_oenb[11]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 937.440 4.000 938.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 742.560 4.000 743.120 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 688.800 1.000 689.360 4.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 43.680 779.000 44.240 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 131.040 1.000 131.600 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 114.240 4.000 114.800 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 991.200 4.000 991.760 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 228.480 779.000 229.040 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 26.880 1076.000 27.440 1079.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 544.320 4.000 544.880 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 231.840 1076.000 232.400 1079.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 537.600 1076.000 538.160 1079.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 258.720 1.000 259.280 4.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 722.400 779.000 722.960 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 50.400 779.000 50.960 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 33.600 1076.000 34.160 1079.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 168.000 1.000 168.560 4.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 571.200 4.000 571.760 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 1034.880 779.000 1035.440 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 769.440 1076.000 770.000 1079.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 947.520 779.000 948.080 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 248.640 1076.000 249.200 1079.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 910.560 779.000 911.120 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 473.760 1.000 474.320 4.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 6.720 1076.000 7.280 1079.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 23.520 1.000 24.080 4.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 6.720 1.000 7.280 4.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1055.040 4.000 1055.600 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 480.480 1.000 481.040 4.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 399.840 4.000 400.400 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 507.360 4.000 507.920 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 265.440 779.000 266.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 188.160 1076.000 188.720 1079.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 588.000 4.000 588.560 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 178.080 1.000 178.640 4.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 409.920 1.000 410.480 4.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 618.240 1076.000 618.800 1079.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 742.560 1.000 743.120 4.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 104.160 4.000 104.720 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 678.720 4.000 679.280 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 6.720 4.000 7.280 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 866.880 4.000 867.440 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 715.680 1.000 716.240 4.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 151.200 1076.000 151.760 1079.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 141.120 779.000 141.680 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 739.200 779.000 739.760 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 500.640 4.000 501.200 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 631.680 779.000 632.240 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 705.600 1.000 706.160 4.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 672.000 1076.000 672.560 1079.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 248.640 779.000 249.200 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 403.200 1076.000 403.760 1079.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 77.280 779.000 77.840 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 453.600 4.000 454.160 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 114.240 1.000 114.800 4.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 614.880 779.000 615.440 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 221.760 4.000 222.320 ;
    END
  END la_oenb[63]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 759.360 779.000 759.920 ;
    END
  END la_oenb[6]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 231.840 1.000 232.400 4.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 104.160 779.000 104.720 ;
    END
  END la_oenb[8]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 114.240 1076.000 114.800 1079.000 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 645.120 1076.000 645.680 1079.000 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 866.880 779.000 867.440 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 80.640 1076.000 81.200 1079.000 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 598.080 4.000 598.640 ;
    END
  END user_irq[2]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 1062.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 1062.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 1062.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 1062.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 1062.620 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 1062.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 1062.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 1062.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 1062.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 1062.620 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 309.120 779.000 309.680 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 16.800 1076.000 17.360 1079.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 470.400 779.000 470.960 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 463.680 1076.000 464.240 1079.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 268.800 1076.000 269.360 1079.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 534.240 4.000 534.800 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 77.280 1.000 77.840 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 517.440 1.000 518.000 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 87.360 4.000 87.920 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 776.160 779.000 776.720 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 588.000 1.000 588.560 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 517.440 4.000 518.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 443.520 779.000 444.080 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 114.240 779.000 114.800 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 60.480 4.000 61.040 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 715.680 1076.000 716.240 1079.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 527.520 1.000 528.080 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 749.280 1.000 749.840 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 362.880 779.000 363.440 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1034.880 4.000 1035.440 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 157.920 4.000 158.480 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 97.440 1.000 98.000 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 161.280 1076.000 161.840 1079.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 695.520 779.000 696.080 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 1044.960 779.000 1045.520 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 366.240 1.000 366.800 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 366.240 4.000 366.800 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 544.320 779.000 544.880 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 722.400 1.000 722.960 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 564.480 1076.000 565.040 1079.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 695.520 1.000 696.080 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 231.840 4.000 232.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 43.680 1.000 44.240 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 151.200 779.000 151.760 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 399.840 779.000 400.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 141.120 1076.000 141.680 1079.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 964.320 779.000 964.880 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 715.680 4.000 716.240 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 786.240 4.000 786.800 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 749.280 4.000 749.840 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 33.600 1.000 34.160 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 194.880 4.000 195.440 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 641.760 779.000 642.320 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 534.240 1.000 534.800 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 483.840 1076.000 484.400 1079.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 705.600 1076.000 706.160 1079.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 981.120 4.000 981.680 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 141.120 1.000 141.680 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 436.800 4.000 437.360 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 732.480 1076.000 733.040 1079.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 554.400 4.000 554.960 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 883.680 779.000 884.240 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 453.600 779.000 454.160 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 641.760 1.000 642.320 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 624.960 1076.000 625.520 1079.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 70.560 1076.000 71.120 1079.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 292.320 1.000 292.880 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 712.320 779.000 712.880 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 759.360 1.000 759.920 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 426.720 779.000 427.280 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 490.560 4.000 491.120 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 184.800 779.000 185.360 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 151.200 1.000 151.760 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 463.680 1.000 464.240 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 551.040 779.000 551.600 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 581.280 1076.000 581.840 1079.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 981.120 779.000 981.680 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 201.600 779.000 202.160 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 184.800 4.000 185.360 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 685.440 779.000 686.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 16.800 1.000 17.360 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 1008.000 779.000 1008.560 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 544.320 1076.000 544.880 1079.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 255.360 779.000 255.920 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 517.440 1076.000 518.000 1079.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 258.720 4.000 259.280 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 292.320 4.000 292.880 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 624.960 1.000 625.520 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1.000 0.560 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 732.480 1.000 733.040 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 446.880 4.000 447.440 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 803.040 4.000 803.600 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 107.520 1076.000 108.080 1079.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 302.400 4.000 302.960 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 194.880 1.000 195.440 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 70.560 1.000 71.120 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 329.280 1076.000 329.840 1079.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 1076.000 124.880 1079.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 507.360 1.000 507.920 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 490.560 1076.000 491.120 1079.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 409.920 779.000 410.480 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 608.160 4.000 608.720 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 873.600 779.000 874.160 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 204.960 1.000 205.520 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 356.160 1.000 356.720 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 77.280 4.000 77.840 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 840.000 779.000 840.560 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 561.120 1.000 561.680 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 456.960 1076.000 457.520 1079.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 446.880 1076.000 447.440 1079.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 856.800 4.000 857.360 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1028.160 4.000 1028.720 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 668.640 1.000 669.200 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 204.960 4.000 205.520 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 769.440 4.000 770.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 776.000 604.800 779.000 605.360 ;
    END
  END wbs_we_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 8.550 776.630 1063.290 ;
      LAYER Metal2 ;
        RECT 0.860 1075.700 6.420 1076.000 ;
        RECT 7.580 1075.700 16.500 1076.000 ;
        RECT 17.660 1075.700 26.580 1076.000 ;
        RECT 27.740 1075.700 33.300 1076.000 ;
        RECT 34.460 1075.700 43.380 1076.000 ;
        RECT 44.540 1075.700 53.460 1076.000 ;
        RECT 54.620 1075.700 60.180 1076.000 ;
        RECT 61.340 1075.700 70.260 1076.000 ;
        RECT 71.420 1075.700 80.340 1076.000 ;
        RECT 81.500 1075.700 87.060 1076.000 ;
        RECT 88.220 1075.700 97.140 1076.000 ;
        RECT 98.300 1075.700 107.220 1076.000 ;
        RECT 108.380 1075.700 113.940 1076.000 ;
        RECT 115.100 1075.700 124.020 1076.000 ;
        RECT 125.180 1075.700 134.100 1076.000 ;
        RECT 135.260 1075.700 140.820 1076.000 ;
        RECT 141.980 1075.700 150.900 1076.000 ;
        RECT 152.060 1075.700 160.980 1076.000 ;
        RECT 162.140 1075.700 167.700 1076.000 ;
        RECT 168.860 1075.700 177.780 1076.000 ;
        RECT 178.940 1075.700 187.860 1076.000 ;
        RECT 189.020 1075.700 194.580 1076.000 ;
        RECT 195.740 1075.700 204.660 1076.000 ;
        RECT 205.820 1075.700 214.740 1076.000 ;
        RECT 215.900 1075.700 221.460 1076.000 ;
        RECT 222.620 1075.700 231.540 1076.000 ;
        RECT 232.700 1075.700 241.620 1076.000 ;
        RECT 242.780 1075.700 248.340 1076.000 ;
        RECT 249.500 1075.700 258.420 1076.000 ;
        RECT 259.580 1075.700 268.500 1076.000 ;
        RECT 269.660 1075.700 275.220 1076.000 ;
        RECT 276.380 1075.700 285.300 1076.000 ;
        RECT 286.460 1075.700 295.380 1076.000 ;
        RECT 296.540 1075.700 302.100 1076.000 ;
        RECT 303.260 1075.700 312.180 1076.000 ;
        RECT 313.340 1075.700 322.260 1076.000 ;
        RECT 323.420 1075.700 328.980 1076.000 ;
        RECT 330.140 1075.700 339.060 1076.000 ;
        RECT 340.220 1075.700 349.140 1076.000 ;
        RECT 350.300 1075.700 355.860 1076.000 ;
        RECT 357.020 1075.700 365.940 1076.000 ;
        RECT 367.100 1075.700 376.020 1076.000 ;
        RECT 377.180 1075.700 382.740 1076.000 ;
        RECT 383.900 1075.700 392.820 1076.000 ;
        RECT 393.980 1075.700 402.900 1076.000 ;
        RECT 404.060 1075.700 409.620 1076.000 ;
        RECT 410.780 1075.700 419.700 1076.000 ;
        RECT 420.860 1075.700 429.780 1076.000 ;
        RECT 430.940 1075.700 436.500 1076.000 ;
        RECT 437.660 1075.700 446.580 1076.000 ;
        RECT 447.740 1075.700 456.660 1076.000 ;
        RECT 457.820 1075.700 463.380 1076.000 ;
        RECT 464.540 1075.700 473.460 1076.000 ;
        RECT 474.620 1075.700 483.540 1076.000 ;
        RECT 484.700 1075.700 490.260 1076.000 ;
        RECT 491.420 1075.700 500.340 1076.000 ;
        RECT 501.500 1075.700 510.420 1076.000 ;
        RECT 511.580 1075.700 517.140 1076.000 ;
        RECT 518.300 1075.700 527.220 1076.000 ;
        RECT 528.380 1075.700 537.300 1076.000 ;
        RECT 538.460 1075.700 544.020 1076.000 ;
        RECT 545.180 1075.700 554.100 1076.000 ;
        RECT 555.260 1075.700 564.180 1076.000 ;
        RECT 565.340 1075.700 570.900 1076.000 ;
        RECT 572.060 1075.700 580.980 1076.000 ;
        RECT 582.140 1075.700 591.060 1076.000 ;
        RECT 592.220 1075.700 597.780 1076.000 ;
        RECT 598.940 1075.700 607.860 1076.000 ;
        RECT 609.020 1075.700 617.940 1076.000 ;
        RECT 619.100 1075.700 624.660 1076.000 ;
        RECT 625.820 1075.700 634.740 1076.000 ;
        RECT 635.900 1075.700 644.820 1076.000 ;
        RECT 645.980 1075.700 651.540 1076.000 ;
        RECT 652.700 1075.700 661.620 1076.000 ;
        RECT 662.780 1075.700 671.700 1076.000 ;
        RECT 672.860 1075.700 678.420 1076.000 ;
        RECT 679.580 1075.700 688.500 1076.000 ;
        RECT 689.660 1075.700 698.580 1076.000 ;
        RECT 699.740 1075.700 705.300 1076.000 ;
        RECT 706.460 1075.700 715.380 1076.000 ;
        RECT 716.540 1075.700 725.460 1076.000 ;
        RECT 726.620 1075.700 732.180 1076.000 ;
        RECT 733.340 1075.700 742.260 1076.000 ;
        RECT 743.420 1075.700 752.340 1076.000 ;
        RECT 753.500 1075.700 759.060 1076.000 ;
        RECT 760.220 1075.700 769.140 1076.000 ;
        RECT 770.300 1075.700 775.860 1076.000 ;
        RECT 0.140 4.300 776.580 1075.700 ;
        RECT 0.860 4.000 6.420 4.300 ;
        RECT 7.580 4.000 16.500 4.300 ;
        RECT 17.660 4.000 23.220 4.300 ;
        RECT 24.380 4.000 33.300 4.300 ;
        RECT 34.460 4.000 43.380 4.300 ;
        RECT 44.540 4.000 50.100 4.300 ;
        RECT 51.260 4.000 60.180 4.300 ;
        RECT 61.340 4.000 70.260 4.300 ;
        RECT 71.420 4.000 76.980 4.300 ;
        RECT 78.140 4.000 87.060 4.300 ;
        RECT 88.220 4.000 97.140 4.300 ;
        RECT 98.300 4.000 103.860 4.300 ;
        RECT 105.020 4.000 113.940 4.300 ;
        RECT 115.100 4.000 124.020 4.300 ;
        RECT 125.180 4.000 130.740 4.300 ;
        RECT 131.900 4.000 140.820 4.300 ;
        RECT 141.980 4.000 150.900 4.300 ;
        RECT 152.060 4.000 157.620 4.300 ;
        RECT 158.780 4.000 167.700 4.300 ;
        RECT 168.860 4.000 177.780 4.300 ;
        RECT 178.940 4.000 184.500 4.300 ;
        RECT 185.660 4.000 194.580 4.300 ;
        RECT 195.740 4.000 204.660 4.300 ;
        RECT 205.820 4.000 211.380 4.300 ;
        RECT 212.540 4.000 221.460 4.300 ;
        RECT 222.620 4.000 231.540 4.300 ;
        RECT 232.700 4.000 238.260 4.300 ;
        RECT 239.420 4.000 248.340 4.300 ;
        RECT 249.500 4.000 258.420 4.300 ;
        RECT 259.580 4.000 265.140 4.300 ;
        RECT 266.300 4.000 275.220 4.300 ;
        RECT 276.380 4.000 285.300 4.300 ;
        RECT 286.460 4.000 292.020 4.300 ;
        RECT 293.180 4.000 302.100 4.300 ;
        RECT 303.260 4.000 312.180 4.300 ;
        RECT 313.340 4.000 318.900 4.300 ;
        RECT 320.060 4.000 328.980 4.300 ;
        RECT 330.140 4.000 339.060 4.300 ;
        RECT 340.220 4.000 345.780 4.300 ;
        RECT 346.940 4.000 355.860 4.300 ;
        RECT 357.020 4.000 365.940 4.300 ;
        RECT 367.100 4.000 372.660 4.300 ;
        RECT 373.820 4.000 382.740 4.300 ;
        RECT 383.900 4.000 392.820 4.300 ;
        RECT 393.980 4.000 399.540 4.300 ;
        RECT 400.700 4.000 409.620 4.300 ;
        RECT 410.780 4.000 419.700 4.300 ;
        RECT 420.860 4.000 426.420 4.300 ;
        RECT 427.580 4.000 436.500 4.300 ;
        RECT 437.660 4.000 446.580 4.300 ;
        RECT 447.740 4.000 453.300 4.300 ;
        RECT 454.460 4.000 463.380 4.300 ;
        RECT 464.540 4.000 473.460 4.300 ;
        RECT 474.620 4.000 480.180 4.300 ;
        RECT 481.340 4.000 490.260 4.300 ;
        RECT 491.420 4.000 500.340 4.300 ;
        RECT 501.500 4.000 507.060 4.300 ;
        RECT 508.220 4.000 517.140 4.300 ;
        RECT 518.300 4.000 527.220 4.300 ;
        RECT 528.380 4.000 533.940 4.300 ;
        RECT 535.100 4.000 544.020 4.300 ;
        RECT 545.180 4.000 554.100 4.300 ;
        RECT 555.260 4.000 560.820 4.300 ;
        RECT 561.980 4.000 570.900 4.300 ;
        RECT 572.060 4.000 580.980 4.300 ;
        RECT 582.140 4.000 587.700 4.300 ;
        RECT 588.860 4.000 597.780 4.300 ;
        RECT 598.940 4.000 607.860 4.300 ;
        RECT 609.020 4.000 614.580 4.300 ;
        RECT 615.740 4.000 624.660 4.300 ;
        RECT 625.820 4.000 634.740 4.300 ;
        RECT 635.900 4.000 641.460 4.300 ;
        RECT 642.620 4.000 651.540 4.300 ;
        RECT 652.700 4.000 661.620 4.300 ;
        RECT 662.780 4.000 668.340 4.300 ;
        RECT 669.500 4.000 678.420 4.300 ;
        RECT 679.580 4.000 688.500 4.300 ;
        RECT 689.660 4.000 695.220 4.300 ;
        RECT 696.380 4.000 705.300 4.300 ;
        RECT 706.460 4.000 715.380 4.300 ;
        RECT 716.540 4.000 722.100 4.300 ;
        RECT 723.260 4.000 732.180 4.300 ;
        RECT 733.340 4.000 742.260 4.300 ;
        RECT 743.420 4.000 748.980 4.300 ;
        RECT 750.140 4.000 759.060 4.300 ;
        RECT 760.220 4.000 769.140 4.300 ;
        RECT 770.300 4.000 775.860 4.300 ;
      LAYER Metal3 ;
        RECT 0.090 1071.540 0.700 1072.260 ;
        RECT 4.300 1071.540 775.700 1072.260 ;
        RECT 0.090 1062.620 776.580 1071.540 ;
        RECT 0.090 1061.460 0.700 1062.620 ;
        RECT 4.300 1061.460 775.700 1062.620 ;
        RECT 0.090 1055.900 776.580 1061.460 ;
        RECT 0.090 1054.740 0.700 1055.900 ;
        RECT 4.300 1054.740 775.700 1055.900 ;
        RECT 0.090 1045.820 776.580 1054.740 ;
        RECT 0.090 1044.660 0.700 1045.820 ;
        RECT 4.300 1044.660 775.700 1045.820 ;
        RECT 0.090 1035.740 776.580 1044.660 ;
        RECT 0.090 1034.580 0.700 1035.740 ;
        RECT 4.300 1034.580 775.700 1035.740 ;
        RECT 0.090 1029.020 776.580 1034.580 ;
        RECT 0.090 1027.860 0.700 1029.020 ;
        RECT 4.300 1027.860 775.700 1029.020 ;
        RECT 0.090 1018.940 776.580 1027.860 ;
        RECT 0.090 1017.780 0.700 1018.940 ;
        RECT 4.300 1017.780 775.700 1018.940 ;
        RECT 0.090 1008.860 776.580 1017.780 ;
        RECT 0.090 1007.700 0.700 1008.860 ;
        RECT 4.300 1007.700 775.700 1008.860 ;
        RECT 0.090 1002.140 776.580 1007.700 ;
        RECT 0.090 1000.980 0.700 1002.140 ;
        RECT 4.300 1000.980 775.700 1002.140 ;
        RECT 0.090 992.060 776.580 1000.980 ;
        RECT 0.090 990.900 0.700 992.060 ;
        RECT 4.300 990.900 775.700 992.060 ;
        RECT 0.090 981.980 776.580 990.900 ;
        RECT 0.090 980.820 0.700 981.980 ;
        RECT 4.300 980.820 775.700 981.980 ;
        RECT 0.090 975.260 776.580 980.820 ;
        RECT 0.090 974.100 0.700 975.260 ;
        RECT 4.300 974.100 775.700 975.260 ;
        RECT 0.090 965.180 776.580 974.100 ;
        RECT 0.090 964.020 0.700 965.180 ;
        RECT 4.300 964.020 775.700 965.180 ;
        RECT 0.090 955.100 776.580 964.020 ;
        RECT 0.090 953.940 0.700 955.100 ;
        RECT 4.300 953.940 775.700 955.100 ;
        RECT 0.090 948.380 776.580 953.940 ;
        RECT 0.090 947.220 0.700 948.380 ;
        RECT 4.300 947.220 775.700 948.380 ;
        RECT 0.090 938.300 776.580 947.220 ;
        RECT 0.090 937.140 0.700 938.300 ;
        RECT 4.300 937.140 775.700 938.300 ;
        RECT 0.090 928.220 776.580 937.140 ;
        RECT 0.090 927.060 0.700 928.220 ;
        RECT 4.300 927.060 775.700 928.220 ;
        RECT 0.090 921.500 776.580 927.060 ;
        RECT 0.090 920.340 0.700 921.500 ;
        RECT 4.300 920.340 775.700 921.500 ;
        RECT 0.090 911.420 776.580 920.340 ;
        RECT 0.090 910.260 0.700 911.420 ;
        RECT 4.300 910.260 775.700 911.420 ;
        RECT 0.090 904.700 776.580 910.260 ;
        RECT 0.090 903.540 0.700 904.700 ;
        RECT 4.300 903.540 776.580 904.700 ;
        RECT 0.090 901.340 776.580 903.540 ;
        RECT 0.090 900.180 775.700 901.340 ;
        RECT 0.090 894.620 776.580 900.180 ;
        RECT 0.090 893.460 0.700 894.620 ;
        RECT 4.300 893.460 775.700 894.620 ;
        RECT 0.090 884.540 776.580 893.460 ;
        RECT 0.090 883.380 0.700 884.540 ;
        RECT 4.300 883.380 775.700 884.540 ;
        RECT 0.090 877.820 776.580 883.380 ;
        RECT 0.090 876.660 0.700 877.820 ;
        RECT 4.300 876.660 776.580 877.820 ;
        RECT 0.090 874.460 776.580 876.660 ;
        RECT 0.090 873.300 775.700 874.460 ;
        RECT 0.090 867.740 776.580 873.300 ;
        RECT 0.090 866.580 0.700 867.740 ;
        RECT 4.300 866.580 775.700 867.740 ;
        RECT 0.090 857.660 776.580 866.580 ;
        RECT 0.090 856.500 0.700 857.660 ;
        RECT 4.300 856.500 775.700 857.660 ;
        RECT 0.090 850.940 776.580 856.500 ;
        RECT 0.090 849.780 0.700 850.940 ;
        RECT 4.300 849.780 776.580 850.940 ;
        RECT 0.090 847.580 776.580 849.780 ;
        RECT 0.090 846.420 775.700 847.580 ;
        RECT 0.090 840.860 776.580 846.420 ;
        RECT 0.090 839.700 0.700 840.860 ;
        RECT 4.300 839.700 775.700 840.860 ;
        RECT 0.090 830.780 776.580 839.700 ;
        RECT 0.090 829.620 0.700 830.780 ;
        RECT 4.300 829.620 775.700 830.780 ;
        RECT 0.090 824.060 776.580 829.620 ;
        RECT 0.090 822.900 0.700 824.060 ;
        RECT 4.300 822.900 776.580 824.060 ;
        RECT 0.090 820.700 776.580 822.900 ;
        RECT 0.090 819.540 775.700 820.700 ;
        RECT 0.090 813.980 776.580 819.540 ;
        RECT 0.090 812.820 0.700 813.980 ;
        RECT 4.300 812.820 775.700 813.980 ;
        RECT 0.090 803.900 776.580 812.820 ;
        RECT 0.090 802.740 0.700 803.900 ;
        RECT 4.300 802.740 775.700 803.900 ;
        RECT 0.090 797.180 776.580 802.740 ;
        RECT 0.090 796.020 0.700 797.180 ;
        RECT 4.300 796.020 776.580 797.180 ;
        RECT 0.090 793.820 776.580 796.020 ;
        RECT 0.090 792.660 775.700 793.820 ;
        RECT 0.090 787.100 776.580 792.660 ;
        RECT 0.090 785.940 0.700 787.100 ;
        RECT 4.300 785.940 775.700 787.100 ;
        RECT 0.090 777.020 776.580 785.940 ;
        RECT 0.090 775.860 0.700 777.020 ;
        RECT 4.300 775.860 775.700 777.020 ;
        RECT 0.090 770.300 776.580 775.860 ;
        RECT 0.090 769.140 0.700 770.300 ;
        RECT 4.300 769.140 776.580 770.300 ;
        RECT 0.090 766.940 776.580 769.140 ;
        RECT 0.090 765.780 775.700 766.940 ;
        RECT 0.090 760.220 776.580 765.780 ;
        RECT 0.090 759.060 0.700 760.220 ;
        RECT 4.300 759.060 775.700 760.220 ;
        RECT 0.090 750.140 776.580 759.060 ;
        RECT 0.090 748.980 0.700 750.140 ;
        RECT 4.300 748.980 775.700 750.140 ;
        RECT 0.090 743.420 776.580 748.980 ;
        RECT 0.090 742.260 0.700 743.420 ;
        RECT 4.300 742.260 776.580 743.420 ;
        RECT 0.090 740.060 776.580 742.260 ;
        RECT 0.090 738.900 775.700 740.060 ;
        RECT 0.090 733.340 776.580 738.900 ;
        RECT 0.090 732.180 0.700 733.340 ;
        RECT 4.300 732.180 775.700 733.340 ;
        RECT 0.090 723.260 776.580 732.180 ;
        RECT 0.090 722.100 0.700 723.260 ;
        RECT 4.300 722.100 775.700 723.260 ;
        RECT 0.090 716.540 776.580 722.100 ;
        RECT 0.090 715.380 0.700 716.540 ;
        RECT 4.300 715.380 776.580 716.540 ;
        RECT 0.090 713.180 776.580 715.380 ;
        RECT 0.090 712.020 775.700 713.180 ;
        RECT 0.090 706.460 776.580 712.020 ;
        RECT 0.090 705.300 0.700 706.460 ;
        RECT 4.300 705.300 775.700 706.460 ;
        RECT 0.090 696.380 776.580 705.300 ;
        RECT 0.090 695.220 0.700 696.380 ;
        RECT 4.300 695.220 775.700 696.380 ;
        RECT 0.090 689.660 776.580 695.220 ;
        RECT 0.090 688.500 0.700 689.660 ;
        RECT 4.300 688.500 776.580 689.660 ;
        RECT 0.090 686.300 776.580 688.500 ;
        RECT 0.090 685.140 775.700 686.300 ;
        RECT 0.090 679.580 776.580 685.140 ;
        RECT 0.090 678.420 0.700 679.580 ;
        RECT 4.300 678.420 775.700 679.580 ;
        RECT 0.090 669.500 776.580 678.420 ;
        RECT 0.090 668.340 0.700 669.500 ;
        RECT 4.300 668.340 775.700 669.500 ;
        RECT 0.090 662.780 776.580 668.340 ;
        RECT 0.090 661.620 0.700 662.780 ;
        RECT 4.300 661.620 776.580 662.780 ;
        RECT 0.090 659.420 776.580 661.620 ;
        RECT 0.090 658.260 775.700 659.420 ;
        RECT 0.090 652.700 776.580 658.260 ;
        RECT 0.090 651.540 0.700 652.700 ;
        RECT 4.300 651.540 775.700 652.700 ;
        RECT 0.090 642.620 776.580 651.540 ;
        RECT 0.090 641.460 0.700 642.620 ;
        RECT 4.300 641.460 775.700 642.620 ;
        RECT 0.090 635.900 776.580 641.460 ;
        RECT 0.090 634.740 0.700 635.900 ;
        RECT 4.300 634.740 776.580 635.900 ;
        RECT 0.090 632.540 776.580 634.740 ;
        RECT 0.090 631.380 775.700 632.540 ;
        RECT 0.090 625.820 776.580 631.380 ;
        RECT 0.090 624.660 0.700 625.820 ;
        RECT 4.300 624.660 775.700 625.820 ;
        RECT 0.090 615.740 776.580 624.660 ;
        RECT 0.090 614.580 0.700 615.740 ;
        RECT 4.300 614.580 775.700 615.740 ;
        RECT 0.090 609.020 776.580 614.580 ;
        RECT 0.090 607.860 0.700 609.020 ;
        RECT 4.300 607.860 776.580 609.020 ;
        RECT 0.090 605.660 776.580 607.860 ;
        RECT 0.090 604.500 775.700 605.660 ;
        RECT 0.090 598.940 776.580 604.500 ;
        RECT 0.090 597.780 0.700 598.940 ;
        RECT 4.300 597.780 775.700 598.940 ;
        RECT 0.090 588.860 776.580 597.780 ;
        RECT 0.090 587.700 0.700 588.860 ;
        RECT 4.300 587.700 775.700 588.860 ;
        RECT 0.090 582.140 776.580 587.700 ;
        RECT 0.090 580.980 0.700 582.140 ;
        RECT 4.300 580.980 776.580 582.140 ;
        RECT 0.090 578.780 776.580 580.980 ;
        RECT 0.090 577.620 775.700 578.780 ;
        RECT 0.090 572.060 776.580 577.620 ;
        RECT 0.090 570.900 0.700 572.060 ;
        RECT 4.300 570.900 775.700 572.060 ;
        RECT 0.090 561.980 776.580 570.900 ;
        RECT 0.090 560.820 0.700 561.980 ;
        RECT 4.300 560.820 775.700 561.980 ;
        RECT 0.090 555.260 776.580 560.820 ;
        RECT 0.090 554.100 0.700 555.260 ;
        RECT 4.300 554.100 776.580 555.260 ;
        RECT 0.090 551.900 776.580 554.100 ;
        RECT 0.090 550.740 775.700 551.900 ;
        RECT 0.090 545.180 776.580 550.740 ;
        RECT 0.090 544.020 0.700 545.180 ;
        RECT 4.300 544.020 775.700 545.180 ;
        RECT 0.090 535.100 776.580 544.020 ;
        RECT 0.090 533.940 0.700 535.100 ;
        RECT 4.300 533.940 775.700 535.100 ;
        RECT 0.090 528.380 776.580 533.940 ;
        RECT 0.090 527.220 0.700 528.380 ;
        RECT 4.300 527.220 776.580 528.380 ;
        RECT 0.090 525.020 776.580 527.220 ;
        RECT 0.090 523.860 775.700 525.020 ;
        RECT 0.090 518.300 776.580 523.860 ;
        RECT 0.090 517.140 0.700 518.300 ;
        RECT 4.300 517.140 775.700 518.300 ;
        RECT 0.090 508.220 776.580 517.140 ;
        RECT 0.090 507.060 0.700 508.220 ;
        RECT 4.300 507.060 775.700 508.220 ;
        RECT 0.090 501.500 776.580 507.060 ;
        RECT 0.090 500.340 0.700 501.500 ;
        RECT 4.300 500.340 776.580 501.500 ;
        RECT 0.090 498.140 776.580 500.340 ;
        RECT 0.090 496.980 775.700 498.140 ;
        RECT 0.090 491.420 776.580 496.980 ;
        RECT 0.090 490.260 0.700 491.420 ;
        RECT 4.300 490.260 775.700 491.420 ;
        RECT 0.090 481.340 776.580 490.260 ;
        RECT 0.090 480.180 0.700 481.340 ;
        RECT 4.300 480.180 775.700 481.340 ;
        RECT 0.090 474.620 776.580 480.180 ;
        RECT 0.090 473.460 0.700 474.620 ;
        RECT 4.300 473.460 776.580 474.620 ;
        RECT 0.090 471.260 776.580 473.460 ;
        RECT 0.090 470.100 775.700 471.260 ;
        RECT 0.090 464.540 776.580 470.100 ;
        RECT 0.090 463.380 0.700 464.540 ;
        RECT 4.300 463.380 775.700 464.540 ;
        RECT 0.090 454.460 776.580 463.380 ;
        RECT 0.090 453.300 0.700 454.460 ;
        RECT 4.300 453.300 775.700 454.460 ;
        RECT 0.090 447.740 776.580 453.300 ;
        RECT 0.090 446.580 0.700 447.740 ;
        RECT 4.300 446.580 776.580 447.740 ;
        RECT 0.090 444.380 776.580 446.580 ;
        RECT 0.090 443.220 775.700 444.380 ;
        RECT 0.090 437.660 776.580 443.220 ;
        RECT 0.090 436.500 0.700 437.660 ;
        RECT 4.300 436.500 775.700 437.660 ;
        RECT 0.090 427.580 776.580 436.500 ;
        RECT 0.090 426.420 0.700 427.580 ;
        RECT 4.300 426.420 775.700 427.580 ;
        RECT 0.090 420.860 776.580 426.420 ;
        RECT 0.090 419.700 0.700 420.860 ;
        RECT 4.300 419.700 776.580 420.860 ;
        RECT 0.090 417.500 776.580 419.700 ;
        RECT 0.090 416.340 775.700 417.500 ;
        RECT 0.090 410.780 776.580 416.340 ;
        RECT 0.090 409.620 0.700 410.780 ;
        RECT 4.300 409.620 775.700 410.780 ;
        RECT 0.090 400.700 776.580 409.620 ;
        RECT 0.090 399.540 0.700 400.700 ;
        RECT 4.300 399.540 775.700 400.700 ;
        RECT 0.090 393.980 776.580 399.540 ;
        RECT 0.090 392.820 0.700 393.980 ;
        RECT 4.300 392.820 776.580 393.980 ;
        RECT 0.090 390.620 776.580 392.820 ;
        RECT 0.090 389.460 775.700 390.620 ;
        RECT 0.090 383.900 776.580 389.460 ;
        RECT 0.090 382.740 0.700 383.900 ;
        RECT 4.300 382.740 775.700 383.900 ;
        RECT 0.090 373.820 776.580 382.740 ;
        RECT 0.090 372.660 0.700 373.820 ;
        RECT 4.300 372.660 775.700 373.820 ;
        RECT 0.090 367.100 776.580 372.660 ;
        RECT 0.090 365.940 0.700 367.100 ;
        RECT 4.300 365.940 776.580 367.100 ;
        RECT 0.090 363.740 776.580 365.940 ;
        RECT 0.090 362.580 775.700 363.740 ;
        RECT 0.090 357.020 776.580 362.580 ;
        RECT 0.090 355.860 0.700 357.020 ;
        RECT 4.300 355.860 775.700 357.020 ;
        RECT 0.090 346.940 776.580 355.860 ;
        RECT 0.090 345.780 0.700 346.940 ;
        RECT 4.300 345.780 775.700 346.940 ;
        RECT 0.090 340.220 776.580 345.780 ;
        RECT 0.090 339.060 0.700 340.220 ;
        RECT 4.300 339.060 776.580 340.220 ;
        RECT 0.090 336.860 776.580 339.060 ;
        RECT 0.090 335.700 775.700 336.860 ;
        RECT 0.090 330.140 776.580 335.700 ;
        RECT 0.090 328.980 0.700 330.140 ;
        RECT 4.300 328.980 775.700 330.140 ;
        RECT 0.090 320.060 776.580 328.980 ;
        RECT 0.090 318.900 0.700 320.060 ;
        RECT 4.300 318.900 775.700 320.060 ;
        RECT 0.090 313.340 776.580 318.900 ;
        RECT 0.090 312.180 0.700 313.340 ;
        RECT 4.300 312.180 776.580 313.340 ;
        RECT 0.090 309.980 776.580 312.180 ;
        RECT 0.090 308.820 775.700 309.980 ;
        RECT 0.090 303.260 776.580 308.820 ;
        RECT 0.090 302.100 0.700 303.260 ;
        RECT 4.300 302.100 775.700 303.260 ;
        RECT 0.090 293.180 776.580 302.100 ;
        RECT 0.090 292.020 0.700 293.180 ;
        RECT 4.300 292.020 775.700 293.180 ;
        RECT 0.090 286.460 776.580 292.020 ;
        RECT 0.090 285.300 0.700 286.460 ;
        RECT 4.300 285.300 776.580 286.460 ;
        RECT 0.090 283.100 776.580 285.300 ;
        RECT 0.090 281.940 775.700 283.100 ;
        RECT 0.090 276.380 776.580 281.940 ;
        RECT 0.090 275.220 0.700 276.380 ;
        RECT 4.300 275.220 775.700 276.380 ;
        RECT 0.090 266.300 776.580 275.220 ;
        RECT 0.090 265.140 0.700 266.300 ;
        RECT 4.300 265.140 775.700 266.300 ;
        RECT 0.090 259.580 776.580 265.140 ;
        RECT 0.090 258.420 0.700 259.580 ;
        RECT 4.300 258.420 776.580 259.580 ;
        RECT 0.090 256.220 776.580 258.420 ;
        RECT 0.090 255.060 775.700 256.220 ;
        RECT 0.090 249.500 776.580 255.060 ;
        RECT 0.090 248.340 0.700 249.500 ;
        RECT 4.300 248.340 775.700 249.500 ;
        RECT 0.090 239.420 776.580 248.340 ;
        RECT 0.090 238.260 0.700 239.420 ;
        RECT 4.300 238.260 775.700 239.420 ;
        RECT 0.090 232.700 776.580 238.260 ;
        RECT 0.090 231.540 0.700 232.700 ;
        RECT 4.300 231.540 776.580 232.700 ;
        RECT 0.090 229.340 776.580 231.540 ;
        RECT 0.090 228.180 775.700 229.340 ;
        RECT 0.090 222.620 776.580 228.180 ;
        RECT 0.090 221.460 0.700 222.620 ;
        RECT 4.300 221.460 775.700 222.620 ;
        RECT 0.090 212.540 776.580 221.460 ;
        RECT 0.090 211.380 0.700 212.540 ;
        RECT 4.300 211.380 775.700 212.540 ;
        RECT 0.090 205.820 776.580 211.380 ;
        RECT 0.090 204.660 0.700 205.820 ;
        RECT 4.300 204.660 776.580 205.820 ;
        RECT 0.090 202.460 776.580 204.660 ;
        RECT 0.090 201.300 775.700 202.460 ;
        RECT 0.090 195.740 776.580 201.300 ;
        RECT 0.090 194.580 0.700 195.740 ;
        RECT 4.300 194.580 775.700 195.740 ;
        RECT 0.090 185.660 776.580 194.580 ;
        RECT 0.090 184.500 0.700 185.660 ;
        RECT 4.300 184.500 775.700 185.660 ;
        RECT 0.090 178.940 776.580 184.500 ;
        RECT 0.090 177.780 0.700 178.940 ;
        RECT 4.300 177.780 776.580 178.940 ;
        RECT 0.090 175.580 776.580 177.780 ;
        RECT 0.090 174.420 775.700 175.580 ;
        RECT 0.090 168.860 776.580 174.420 ;
        RECT 0.090 167.700 0.700 168.860 ;
        RECT 4.300 167.700 775.700 168.860 ;
        RECT 0.090 158.780 776.580 167.700 ;
        RECT 0.090 157.620 0.700 158.780 ;
        RECT 4.300 157.620 775.700 158.780 ;
        RECT 0.090 152.060 776.580 157.620 ;
        RECT 0.090 150.900 0.700 152.060 ;
        RECT 4.300 150.900 775.700 152.060 ;
        RECT 0.090 141.980 776.580 150.900 ;
        RECT 0.090 140.820 0.700 141.980 ;
        RECT 4.300 140.820 775.700 141.980 ;
        RECT 0.090 131.900 776.580 140.820 ;
        RECT 0.090 130.740 0.700 131.900 ;
        RECT 4.300 130.740 775.700 131.900 ;
        RECT 0.090 125.180 776.580 130.740 ;
        RECT 0.090 124.020 0.700 125.180 ;
        RECT 4.300 124.020 775.700 125.180 ;
        RECT 0.090 115.100 776.580 124.020 ;
        RECT 0.090 113.940 0.700 115.100 ;
        RECT 4.300 113.940 775.700 115.100 ;
        RECT 0.090 105.020 776.580 113.940 ;
        RECT 0.090 103.860 0.700 105.020 ;
        RECT 4.300 103.860 775.700 105.020 ;
        RECT 0.090 98.300 776.580 103.860 ;
        RECT 0.090 97.140 0.700 98.300 ;
        RECT 4.300 97.140 775.700 98.300 ;
        RECT 0.090 88.220 776.580 97.140 ;
        RECT 0.090 87.060 0.700 88.220 ;
        RECT 4.300 87.060 775.700 88.220 ;
        RECT 0.090 78.140 776.580 87.060 ;
        RECT 0.090 76.980 0.700 78.140 ;
        RECT 4.300 76.980 775.700 78.140 ;
        RECT 0.090 71.420 776.580 76.980 ;
        RECT 0.090 70.260 0.700 71.420 ;
        RECT 4.300 70.260 775.700 71.420 ;
        RECT 0.090 61.340 776.580 70.260 ;
        RECT 0.090 60.180 0.700 61.340 ;
        RECT 4.300 60.180 775.700 61.340 ;
        RECT 0.090 51.260 776.580 60.180 ;
        RECT 0.090 50.100 0.700 51.260 ;
        RECT 4.300 50.100 775.700 51.260 ;
        RECT 0.090 44.540 776.580 50.100 ;
        RECT 0.090 43.380 0.700 44.540 ;
        RECT 4.300 43.380 775.700 44.540 ;
        RECT 0.090 34.460 776.580 43.380 ;
        RECT 0.090 33.300 0.700 34.460 ;
        RECT 4.300 33.300 775.700 34.460 ;
        RECT 0.090 24.380 776.580 33.300 ;
        RECT 0.090 23.220 0.700 24.380 ;
        RECT 4.300 23.220 775.700 24.380 ;
        RECT 0.090 17.660 776.580 23.220 ;
        RECT 0.090 16.500 0.700 17.660 ;
        RECT 4.300 16.500 775.700 17.660 ;
        RECT 0.090 7.980 776.580 16.500 ;
      LAYER Metal4 ;
        RECT 16.660 116.010 21.940 924.470 ;
        RECT 24.140 116.010 98.740 924.470 ;
        RECT 100.940 116.010 175.540 924.470 ;
        RECT 177.740 116.010 252.340 924.470 ;
        RECT 254.540 116.010 329.140 924.470 ;
        RECT 331.340 116.010 405.940 924.470 ;
        RECT 408.140 116.010 482.740 924.470 ;
        RECT 484.940 116.010 559.540 924.470 ;
        RECT 561.740 116.010 636.340 924.470 ;
        RECT 638.540 116.010 688.100 924.470 ;
  END
END tiny_user_project
END LIBRARY

