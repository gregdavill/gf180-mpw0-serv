VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tiny_user_project
  CLASS BLOCK ;
  FOREIGN tiny_user_project ;
  ORIGIN 0.000 0.000 ;
  SIZE 690.000 BY 800.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 514.080 4.000 514.640 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 520.800 4.000 521.360 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 255.360 4.000 255.920 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 450.240 4.000 450.800 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 305.760 4.000 306.320 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 262.080 4.000 262.640 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 339.360 796.000 339.920 799.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 201.600 689.000 202.160 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 756.000 689.000 756.560 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 446.880 796.000 447.440 799.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 36.960 689.000 37.520 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 36.960 796.000 37.520 799.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 540.960 796.000 541.520 799.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 520.800 1.000 521.360 4.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 688.800 796.000 689.360 799.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 698.880 689.000 699.440 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 614.880 1.000 615.440 4.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 97.440 1.000 98.000 4.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 621.600 4.000 622.160 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 507.360 4.000 507.920 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 577.920 4.000 578.480 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 463.680 4.000 464.240 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 789.600 689.000 790.160 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 487.200 1.000 487.760 4.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 312.480 4.000 313.040 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 628.320 1.000 628.880 4.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 77.280 4.000 77.840 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 665.280 4.000 665.840 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 611.520 796.000 612.080 799.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 712.320 689.000 712.880 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 618.240 689.000 618.800 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 782.880 689.000 783.440 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 389.760 689.000 390.320 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 141.120 4.000 141.680 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 194.880 689.000 195.440 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 554.400 796.000 554.960 799.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 342.720 4.000 343.280 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 386.400 4.000 386.960 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 574.560 689.000 575.120 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 534.240 689.000 534.800 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 772.800 4.000 773.360 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 456.960 1.000 457.520 4.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 191.520 4.000 192.080 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 678.720 1.000 679.280 4.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 416.640 796.000 417.200 799.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 215.040 1.000 215.600 4.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 70.560 1.000 71.120 4.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 779.520 4.000 780.080 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 208.320 796.000 208.880 799.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 144.480 796.000 145.040 799.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 376.320 796.000 376.880 799.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 635.040 1.000 635.600 4.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 245.280 689.000 245.840 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 668.640 796.000 669.200 799.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 215.040 4.000 215.600 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 107.520 4.000 108.080 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 678.720 4.000 679.280 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 621.600 1.000 622.160 4.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 759.360 4.000 759.920 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 433.440 689.000 434.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 339.360 689.000 339.920 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 10.080 689.000 10.640 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 228.480 4.000 229.040 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 598.080 796.000 598.640 799.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 174.720 689.000 175.280 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 608.160 4.000 608.720 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 725.760 689.000 726.320 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 359.520 796.000 360.080 799.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 352.800 689.000 353.360 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 557.760 4.000 558.320 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 97.440 4.000 98.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 490.560 796.000 491.120 799.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 588.000 4.000 588.560 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 302.400 796.000 302.960 799.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 369.600 4.000 370.160 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 776.160 689.000 776.720 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 67.200 796.000 67.760 799.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 174.720 796.000 175.280 799.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 480.480 1.000 481.040 4.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 675.360 796.000 675.920 799.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 742.560 4.000 743.120 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 551.040 4.000 551.600 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 299.040 1.000 299.600 4.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 675.360 689.000 675.920 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 84.000 1.000 84.560 4.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 3.360 689.000 3.920 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 110.880 796.000 111.440 799.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 47.040 1.000 47.600 4.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 124.320 689.000 124.880 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 493.920 4.000 494.480 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 218.400 689.000 218.960 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 278.880 4.000 279.440 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 651.840 1.000 652.400 4.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 73.920 689.000 74.480 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 312.480 1.000 313.040 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 248.640 1.000 249.200 4.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 467.040 796.000 467.600 799.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 507.360 1.000 507.920 4.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 315.840 689.000 316.400 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 624.960 796.000 625.520 799.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 262.080 1.000 262.640 4.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 409.920 796.000 410.480 799.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 272.160 4.000 272.720 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 493.920 1.000 494.480 4.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 443.520 1.000 444.080 4.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 178.080 1.000 178.640 4.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 33.600 4.000 34.160 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 288.960 796.000 289.520 799.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 342.720 1.000 343.280 4.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 258.720 796.000 259.280 799.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 134.400 4.000 134.960 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 420.000 4.000 420.560 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 544.320 1.000 544.880 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 191.520 1.000 192.080 4.000 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 379.680 4.000 380.240 ;
    END
  END la_data_in[0]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 749.280 689.000 749.840 ;
    END
  END la_data_in[10]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 383.040 689.000 383.600 ;
    END
  END la_data_in[11]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 228.480 1.000 229.040 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 245.280 796.000 245.840 799.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 651.840 4.000 652.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 591.360 689.000 591.920 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 16.800 796.000 17.360 799.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 168.000 689.000 168.560 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 315.840 796.000 316.400 799.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 114.240 4.000 114.800 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 117.600 796.000 118.160 799.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 208.320 689.000 208.880 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 564.480 4.000 565.040 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 329.280 4.000 329.840 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 611.520 689.000 612.080 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 325.920 796.000 326.480 799.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 100.800 796.000 101.360 799.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 403.200 796.000 403.760 799.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 672.000 4.000 672.560 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 702.240 4.000 702.800 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 238.560 689.000 239.120 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 275.520 796.000 276.080 799.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 57.120 4.000 57.680 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 574.560 796.000 575.120 799.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 299.040 4.000 299.600 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 500.640 4.000 501.200 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3.360 796.000 3.920 799.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 658.560 4.000 659.120 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 527.520 1.000 528.080 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 729.120 4.000 729.680 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 336.000 1.000 336.560 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 352.800 796.000 353.360 799.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 460.320 689.000 460.880 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 255.360 1.000 255.920 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 356.160 1.000 356.720 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 248.640 4.000 249.200 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 648.480 796.000 649.040 799.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 60.480 689.000 61.040 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 241.920 1.000 242.480 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 598.080 689.000 598.640 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 463.680 1.000 464.240 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 295.680 796.000 296.240 799.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 231.840 796.000 232.400 799.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 10.080 796.000 10.640 799.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 238.560 796.000 239.120 799.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 349.440 1.000 350.000 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 302.400 689.000 302.960 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 524.160 796.000 524.720 799.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 473.760 796.000 474.320 799.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 198.240 4.000 198.800 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 221.760 4.000 222.320 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 766.080 4.000 766.640 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 272.160 1.000 272.720 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 732.480 689.000 733.040 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 127.680 1.000 128.240 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 547.680 689.000 548.240 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 20.160 4.000 20.720 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 436.800 1.000 437.360 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 137.760 796.000 138.320 799.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 147.840 1.000 148.400 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 325.920 689.000 326.480 ;
    END
  END la_data_in[7]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 13.440 4.000 14.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 618.240 796.000 618.800 799.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 591.360 796.000 591.920 799.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 453.600 689.000 454.160 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 26.880 4.000 27.440 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 537.600 4.000 538.160 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 278.880 1.000 279.440 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 359.520 689.000 360.080 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 635.040 4.000 635.600 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 467.040 689.000 467.600 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 309.120 796.000 309.680 799.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 668.640 689.000 669.200 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 393.120 1.000 393.680 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 403.200 689.000 403.760 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 161.280 689.000 161.840 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 735.840 4.000 736.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 517.440 689.000 518.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 221.760 1.000 222.320 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 336.000 4.000 336.560 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 399.840 1.000 400.400 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 722.400 4.000 722.960 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 396.480 796.000 397.040 799.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 648.480 689.000 649.040 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 322.560 1.000 323.120 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 171.360 4.000 171.920 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 396.480 689.000 397.040 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 87.360 689.000 87.920 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 383.040 796.000 383.600 799.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 188.160 689.000 188.720 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 362.880 1.000 363.440 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 346.080 796.000 346.640 799.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 655.200 689.000 655.760 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 346.080 689.000 346.640 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 67.200 689.000 67.760 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 151.200 689.000 151.760 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 120.960 4.000 121.520 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 30.240 689.000 30.800 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 282.240 689.000 282.800 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 682.080 689.000 682.640 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 40.320 1.000 40.880 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 305.760 1.000 306.320 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 60.480 796.000 61.040 799.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 53.760 796.000 54.320 799.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 527.520 4.000 528.080 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 171.360 1.000 171.920 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 672.000 1.000 672.560 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 366.240 796.000 366.800 799.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 201.600 796.000 202.160 799.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 715.680 4.000 716.240 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 100.800 689.000 101.360 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 708.960 4.000 709.520 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 561.120 689.000 561.680 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 225.120 796.000 225.680 799.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 231.840 689.000 232.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 510.720 796.000 511.280 799.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 567.840 689.000 568.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 285.600 4.000 286.160 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 497.280 689.000 497.840 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 547.680 796.000 548.240 799.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 198.240 1.000 198.800 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 645.120 1.000 645.680 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 110.880 689.000 111.440 ;
    END
  END la_data_out[63]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 268.800 689.000 269.360 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 661.920 796.000 662.480 799.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 40.320 4.000 40.880 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 409.920 689.000 410.480 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 332.640 689.000 333.200 ;
    END
  END la_oenb[0]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 581.280 689.000 581.840 ;
    END
  END la_oenb[10]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 473.760 689.000 474.320 ;
    END
  END la_oenb[11]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 752.640 4.000 753.200 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 594.720 4.000 595.280 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 551.040 1.000 551.600 4.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 658.560 1.000 659.120 4.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 107.520 1.000 108.080 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 90.720 4.000 91.280 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 792.960 4.000 793.520 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 117.600 689.000 118.160 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 87.360 796.000 87.920 799.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 436.800 4.000 437.360 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 252.000 796.000 252.560 799.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 497.280 796.000 497.840 799.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 204.960 1.000 205.520 4.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 510.720 689.000 511.280 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 665.280 1.000 665.840 4.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 94.080 796.000 94.640 799.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 134.400 1.000 134.960 4.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 456.960 4.000 457.520 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 762.720 689.000 763.280 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 682.080 796.000 682.640 799.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 688.800 689.000 689.360 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 268.800 796.000 269.360 799.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 661.920 689.000 662.480 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 379.680 1.000 380.240 4.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 73.920 796.000 74.480 799.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 20.160 1.000 20.720 4.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 6.720 1.000 7.280 4.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 43.680 796.000 44.240 799.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 386.400 1.000 386.960 4.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 322.560 4.000 323.120 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 406.560 4.000 407.120 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 144.480 689.000 145.040 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 218.400 796.000 218.960 799.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 470.400 4.000 470.960 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 141.120 1.000 141.680 4.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 329.280 1.000 329.840 4.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 561.120 796.000 561.680 799.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 594.720 1.000 595.280 4.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 84.000 4.000 84.560 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 544.320 4.000 544.880 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 6.720 4.000 7.280 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 695.520 4.000 696.080 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 571.200 1.000 571.760 4.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 188.160 796.000 188.720 799.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 43.680 689.000 44.240 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 524.160 689.000 524.720 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 399.840 4.000 400.400 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 440.160 689.000 440.720 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 564.480 1.000 565.040 4.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 604.800 796.000 605.360 799.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 131.040 689.000 131.600 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 389.760 796.000 390.320 799.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 685.440 1.000 686.000 4.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 362.880 4.000 363.440 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 1.000 91.280 4.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 426.720 689.000 427.280 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 178.080 4.000 178.640 ;
    END
  END la_oenb[63]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 540.960 689.000 541.520 ;
    END
  END la_oenb[6]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 184.800 1.000 185.360 4.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 16.800 689.000 17.360 ;
    END
  END la_oenb[8]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 161.280 796.000 161.840 799.000 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 581.280 796.000 581.840 799.000 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 624.960 689.000 625.520 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 131.040 796.000 131.600 799.000 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 480.480 4.000 481.040 ;
    END
  END user_irq[2]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 784.300 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 784.300 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 181.440 689.000 182.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 80.640 796.000 81.200 799.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 309.120 689.000 309.680 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 440.160 796.000 440.720 799.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 282.240 796.000 282.800 799.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 430.080 4.000 430.640 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 63.840 1.000 64.400 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 413.280 1.000 413.840 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 70.560 4.000 71.120 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 554.400 689.000 554.960 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 470.400 1.000 470.960 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 413.280 4.000 413.840 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 288.960 689.000 289.520 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 23.520 689.000 24.080 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 47.040 4.000 47.600 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 641.760 796.000 642.320 799.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 420.000 1.000 420.560 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 601.440 1.000 602.000 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 225.120 689.000 225.680 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 30.240 796.000 30.800 799.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 127.680 4.000 128.240 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 77.280 1.000 77.840 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 194.880 796.000 195.440 799.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 490.560 689.000 491.120 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 769.440 689.000 770.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 292.320 1.000 292.880 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 292.320 4.000 292.880 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 366.240 689.000 366.800 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 577.920 1.000 578.480 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 517.440 796.000 518.000 799.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 557.760 1.000 558.320 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 184.800 4.000 185.360 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 33.600 1.000 34.160 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 53.760 689.000 54.320 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 252.000 689.000 252.560 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 181.440 796.000 182.000 799.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 705.600 689.000 706.160 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 571.200 4.000 571.760 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 628.320 4.000 628.880 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 601.440 4.000 602.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 26.880 1.000 27.440 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 154.560 4.000 155.120 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 446.880 689.000 447.440 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 430.080 1.000 430.640 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 453.600 796.000 454.160 799.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 631.680 796.000 632.240 799.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 786.240 4.000 786.800 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 114.240 1.000 114.800 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 349.440 4.000 350.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 655.200 796.000 655.760 799.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 443.520 4.000 444.080 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 641.760 689.000 642.320 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 295.680 689.000 296.240 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 514.080 1.000 514.640 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 567.840 796.000 568.400 799.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 796.000 124.880 799.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 235.200 1.000 235.760 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 504.000 689.000 504.560 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 608.160 1.000 608.720 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 275.520 689.000 276.080 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 393.120 4.000 393.680 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 80.640 689.000 81.200 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 120.960 1.000 121.520 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 372.960 1.000 373.520 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 376.320 689.000 376.880 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 534.240 796.000 534.800 799.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 719.040 689.000 719.600 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 94.080 689.000 94.640 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 147.840 4.000 148.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 483.840 689.000 484.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 13.440 1.000 14.000 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 739.200 689.000 739.760 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 504.000 796.000 504.560 799.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 137.760 689.000 138.320 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 483.840 796.000 484.400 799.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 204.960 4.000 205.520 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 235.200 4.000 235.760 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 500.640 1.000 501.200 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1.000 0.560 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 588.000 1.000 588.560 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 356.160 4.000 356.720 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 645.120 4.000 645.680 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 151.200 796.000 151.760 799.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 241.920 4.000 242.480 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 154.560 1.000 155.120 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 57.120 1.000 57.680 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 332.640 796.000 333.200 799.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 168.000 796.000 168.560 799.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 406.560 1.000 407.120 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 460.320 796.000 460.880 799.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 258.720 689.000 259.280 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 487.200 4.000 487.760 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 631.680 689.000 632.240 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 164.640 1.000 165.200 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 285.600 1.000 286.160 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 63.840 4.000 64.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 604.800 689.000 605.360 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 450.240 1.000 450.800 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 433.440 796.000 434.000 799.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 426.720 796.000 427.280 799.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 685.440 4.000 686.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 23.520 796.000 24.080 799.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 537.600 1.000 538.160 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 164.640 4.000 165.200 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 614.880 4.000 615.440 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 686.000 416.640 689.000 417.200 ;
    END
  END wbs_we_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 8.550 683.200 784.970 ;
      LAYER Metal2 ;
        RECT 0.140 795.700 3.060 796.000 ;
        RECT 4.220 795.700 9.780 796.000 ;
        RECT 10.940 795.700 16.500 796.000 ;
        RECT 17.660 795.700 23.220 796.000 ;
        RECT 24.380 795.700 29.940 796.000 ;
        RECT 31.100 795.700 36.660 796.000 ;
        RECT 37.820 795.700 43.380 796.000 ;
        RECT 44.540 795.700 53.460 796.000 ;
        RECT 54.620 795.700 60.180 796.000 ;
        RECT 61.340 795.700 66.900 796.000 ;
        RECT 68.060 795.700 73.620 796.000 ;
        RECT 74.780 795.700 80.340 796.000 ;
        RECT 81.500 795.700 87.060 796.000 ;
        RECT 88.220 795.700 93.780 796.000 ;
        RECT 94.940 795.700 100.500 796.000 ;
        RECT 101.660 795.700 110.580 796.000 ;
        RECT 111.740 795.700 117.300 796.000 ;
        RECT 118.460 795.700 124.020 796.000 ;
        RECT 125.180 795.700 130.740 796.000 ;
        RECT 131.900 795.700 137.460 796.000 ;
        RECT 138.620 795.700 144.180 796.000 ;
        RECT 145.340 795.700 150.900 796.000 ;
        RECT 152.060 795.700 160.980 796.000 ;
        RECT 162.140 795.700 167.700 796.000 ;
        RECT 168.860 795.700 174.420 796.000 ;
        RECT 175.580 795.700 181.140 796.000 ;
        RECT 182.300 795.700 187.860 796.000 ;
        RECT 189.020 795.700 194.580 796.000 ;
        RECT 195.740 795.700 201.300 796.000 ;
        RECT 202.460 795.700 208.020 796.000 ;
        RECT 209.180 795.700 218.100 796.000 ;
        RECT 219.260 795.700 224.820 796.000 ;
        RECT 225.980 795.700 231.540 796.000 ;
        RECT 232.700 795.700 238.260 796.000 ;
        RECT 239.420 795.700 244.980 796.000 ;
        RECT 246.140 795.700 251.700 796.000 ;
        RECT 252.860 795.700 258.420 796.000 ;
        RECT 259.580 795.700 268.500 796.000 ;
        RECT 269.660 795.700 275.220 796.000 ;
        RECT 276.380 795.700 281.940 796.000 ;
        RECT 283.100 795.700 288.660 796.000 ;
        RECT 289.820 795.700 295.380 796.000 ;
        RECT 296.540 795.700 302.100 796.000 ;
        RECT 303.260 795.700 308.820 796.000 ;
        RECT 309.980 795.700 315.540 796.000 ;
        RECT 316.700 795.700 325.620 796.000 ;
        RECT 326.780 795.700 332.340 796.000 ;
        RECT 333.500 795.700 339.060 796.000 ;
        RECT 340.220 795.700 345.780 796.000 ;
        RECT 346.940 795.700 352.500 796.000 ;
        RECT 353.660 795.700 359.220 796.000 ;
        RECT 360.380 795.700 365.940 796.000 ;
        RECT 367.100 795.700 376.020 796.000 ;
        RECT 377.180 795.700 382.740 796.000 ;
        RECT 383.900 795.700 389.460 796.000 ;
        RECT 390.620 795.700 396.180 796.000 ;
        RECT 397.340 795.700 402.900 796.000 ;
        RECT 404.060 795.700 409.620 796.000 ;
        RECT 410.780 795.700 416.340 796.000 ;
        RECT 417.500 795.700 426.420 796.000 ;
        RECT 427.580 795.700 433.140 796.000 ;
        RECT 434.300 795.700 439.860 796.000 ;
        RECT 441.020 795.700 446.580 796.000 ;
        RECT 447.740 795.700 453.300 796.000 ;
        RECT 454.460 795.700 460.020 796.000 ;
        RECT 461.180 795.700 466.740 796.000 ;
        RECT 467.900 795.700 473.460 796.000 ;
        RECT 474.620 795.700 483.540 796.000 ;
        RECT 484.700 795.700 490.260 796.000 ;
        RECT 491.420 795.700 496.980 796.000 ;
        RECT 498.140 795.700 503.700 796.000 ;
        RECT 504.860 795.700 510.420 796.000 ;
        RECT 511.580 795.700 517.140 796.000 ;
        RECT 518.300 795.700 523.860 796.000 ;
        RECT 525.020 795.700 533.940 796.000 ;
        RECT 535.100 795.700 540.660 796.000 ;
        RECT 541.820 795.700 547.380 796.000 ;
        RECT 548.540 795.700 554.100 796.000 ;
        RECT 555.260 795.700 560.820 796.000 ;
        RECT 561.980 795.700 567.540 796.000 ;
        RECT 568.700 795.700 574.260 796.000 ;
        RECT 575.420 795.700 580.980 796.000 ;
        RECT 582.140 795.700 591.060 796.000 ;
        RECT 592.220 795.700 597.780 796.000 ;
        RECT 598.940 795.700 604.500 796.000 ;
        RECT 605.660 795.700 611.220 796.000 ;
        RECT 612.380 795.700 617.940 796.000 ;
        RECT 619.100 795.700 624.660 796.000 ;
        RECT 625.820 795.700 631.380 796.000 ;
        RECT 632.540 795.700 641.460 796.000 ;
        RECT 642.620 795.700 648.180 796.000 ;
        RECT 649.340 795.700 654.900 796.000 ;
        RECT 656.060 795.700 661.620 796.000 ;
        RECT 662.780 795.700 668.340 796.000 ;
        RECT 669.500 795.700 675.060 796.000 ;
        RECT 676.220 795.700 681.780 796.000 ;
        RECT 682.940 795.700 686.420 796.000 ;
        RECT 0.140 4.300 686.420 795.700 ;
        RECT 0.860 4.000 6.420 4.300 ;
        RECT 7.580 4.000 13.140 4.300 ;
        RECT 14.300 4.000 19.860 4.300 ;
        RECT 21.020 4.000 26.580 4.300 ;
        RECT 27.740 4.000 33.300 4.300 ;
        RECT 34.460 4.000 40.020 4.300 ;
        RECT 41.180 4.000 46.740 4.300 ;
        RECT 47.900 4.000 56.820 4.300 ;
        RECT 57.980 4.000 63.540 4.300 ;
        RECT 64.700 4.000 70.260 4.300 ;
        RECT 71.420 4.000 76.980 4.300 ;
        RECT 78.140 4.000 83.700 4.300 ;
        RECT 84.860 4.000 90.420 4.300 ;
        RECT 91.580 4.000 97.140 4.300 ;
        RECT 98.300 4.000 107.220 4.300 ;
        RECT 108.380 4.000 113.940 4.300 ;
        RECT 115.100 4.000 120.660 4.300 ;
        RECT 121.820 4.000 127.380 4.300 ;
        RECT 128.540 4.000 134.100 4.300 ;
        RECT 135.260 4.000 140.820 4.300 ;
        RECT 141.980 4.000 147.540 4.300 ;
        RECT 148.700 4.000 154.260 4.300 ;
        RECT 155.420 4.000 164.340 4.300 ;
        RECT 165.500 4.000 171.060 4.300 ;
        RECT 172.220 4.000 177.780 4.300 ;
        RECT 178.940 4.000 184.500 4.300 ;
        RECT 185.660 4.000 191.220 4.300 ;
        RECT 192.380 4.000 197.940 4.300 ;
        RECT 199.100 4.000 204.660 4.300 ;
        RECT 205.820 4.000 214.740 4.300 ;
        RECT 215.900 4.000 221.460 4.300 ;
        RECT 222.620 4.000 228.180 4.300 ;
        RECT 229.340 4.000 234.900 4.300 ;
        RECT 236.060 4.000 241.620 4.300 ;
        RECT 242.780 4.000 248.340 4.300 ;
        RECT 249.500 4.000 255.060 4.300 ;
        RECT 256.220 4.000 261.780 4.300 ;
        RECT 262.940 4.000 271.860 4.300 ;
        RECT 273.020 4.000 278.580 4.300 ;
        RECT 279.740 4.000 285.300 4.300 ;
        RECT 286.460 4.000 292.020 4.300 ;
        RECT 293.180 4.000 298.740 4.300 ;
        RECT 299.900 4.000 305.460 4.300 ;
        RECT 306.620 4.000 312.180 4.300 ;
        RECT 313.340 4.000 322.260 4.300 ;
        RECT 323.420 4.000 328.980 4.300 ;
        RECT 330.140 4.000 335.700 4.300 ;
        RECT 336.860 4.000 342.420 4.300 ;
        RECT 343.580 4.000 349.140 4.300 ;
        RECT 350.300 4.000 355.860 4.300 ;
        RECT 357.020 4.000 362.580 4.300 ;
        RECT 363.740 4.000 372.660 4.300 ;
        RECT 373.820 4.000 379.380 4.300 ;
        RECT 380.540 4.000 386.100 4.300 ;
        RECT 387.260 4.000 392.820 4.300 ;
        RECT 393.980 4.000 399.540 4.300 ;
        RECT 400.700 4.000 406.260 4.300 ;
        RECT 407.420 4.000 412.980 4.300 ;
        RECT 414.140 4.000 419.700 4.300 ;
        RECT 420.860 4.000 429.780 4.300 ;
        RECT 430.940 4.000 436.500 4.300 ;
        RECT 437.660 4.000 443.220 4.300 ;
        RECT 444.380 4.000 449.940 4.300 ;
        RECT 451.100 4.000 456.660 4.300 ;
        RECT 457.820 4.000 463.380 4.300 ;
        RECT 464.540 4.000 470.100 4.300 ;
        RECT 471.260 4.000 480.180 4.300 ;
        RECT 481.340 4.000 486.900 4.300 ;
        RECT 488.060 4.000 493.620 4.300 ;
        RECT 494.780 4.000 500.340 4.300 ;
        RECT 501.500 4.000 507.060 4.300 ;
        RECT 508.220 4.000 513.780 4.300 ;
        RECT 514.940 4.000 520.500 4.300 ;
        RECT 521.660 4.000 527.220 4.300 ;
        RECT 528.380 4.000 537.300 4.300 ;
        RECT 538.460 4.000 544.020 4.300 ;
        RECT 545.180 4.000 550.740 4.300 ;
        RECT 551.900 4.000 557.460 4.300 ;
        RECT 558.620 4.000 564.180 4.300 ;
        RECT 565.340 4.000 570.900 4.300 ;
        RECT 572.060 4.000 577.620 4.300 ;
        RECT 578.780 4.000 587.700 4.300 ;
        RECT 588.860 4.000 594.420 4.300 ;
        RECT 595.580 4.000 601.140 4.300 ;
        RECT 602.300 4.000 607.860 4.300 ;
        RECT 609.020 4.000 614.580 4.300 ;
        RECT 615.740 4.000 621.300 4.300 ;
        RECT 622.460 4.000 628.020 4.300 ;
        RECT 629.180 4.000 634.740 4.300 ;
        RECT 635.900 4.000 644.820 4.300 ;
        RECT 645.980 4.000 651.540 4.300 ;
        RECT 652.700 4.000 658.260 4.300 ;
        RECT 659.420 4.000 664.980 4.300 ;
        RECT 666.140 4.000 671.700 4.300 ;
        RECT 672.860 4.000 678.420 4.300 ;
        RECT 679.580 4.000 685.140 4.300 ;
        RECT 686.300 4.000 686.420 4.300 ;
      LAYER Metal3 ;
        RECT 0.090 783.740 689.780 784.140 ;
        RECT 0.090 782.580 685.700 783.740 ;
        RECT 689.300 782.580 689.780 783.740 ;
        RECT 0.090 780.380 689.780 782.580 ;
        RECT 0.090 779.220 0.700 780.380 ;
        RECT 4.300 779.220 689.780 780.380 ;
        RECT 0.090 777.020 689.780 779.220 ;
        RECT 0.090 775.860 685.700 777.020 ;
        RECT 689.300 775.860 689.780 777.020 ;
        RECT 0.090 773.660 689.780 775.860 ;
        RECT 0.090 772.500 0.700 773.660 ;
        RECT 4.300 772.500 689.780 773.660 ;
        RECT 0.090 770.300 689.780 772.500 ;
        RECT 0.090 769.140 685.700 770.300 ;
        RECT 689.300 769.140 689.780 770.300 ;
        RECT 0.090 766.940 689.780 769.140 ;
        RECT 0.090 765.780 0.700 766.940 ;
        RECT 4.300 765.780 689.780 766.940 ;
        RECT 0.090 763.580 689.780 765.780 ;
        RECT 0.090 762.420 685.700 763.580 ;
        RECT 689.300 762.420 689.780 763.580 ;
        RECT 0.090 760.220 689.780 762.420 ;
        RECT 0.090 759.060 0.700 760.220 ;
        RECT 4.300 759.060 689.780 760.220 ;
        RECT 0.090 756.860 689.780 759.060 ;
        RECT 0.090 755.700 685.700 756.860 ;
        RECT 689.300 755.700 689.780 756.860 ;
        RECT 0.090 753.500 689.780 755.700 ;
        RECT 0.090 752.340 0.700 753.500 ;
        RECT 4.300 752.340 689.780 753.500 ;
        RECT 0.090 750.140 689.780 752.340 ;
        RECT 0.090 748.980 685.700 750.140 ;
        RECT 689.300 748.980 689.780 750.140 ;
        RECT 0.090 743.420 689.780 748.980 ;
        RECT 0.090 742.260 0.700 743.420 ;
        RECT 4.300 742.260 689.780 743.420 ;
        RECT 0.090 740.060 689.780 742.260 ;
        RECT 0.090 738.900 685.700 740.060 ;
        RECT 689.300 738.900 689.780 740.060 ;
        RECT 0.090 736.700 689.780 738.900 ;
        RECT 0.090 735.540 0.700 736.700 ;
        RECT 4.300 735.540 689.780 736.700 ;
        RECT 0.090 733.340 689.780 735.540 ;
        RECT 0.090 732.180 685.700 733.340 ;
        RECT 689.300 732.180 689.780 733.340 ;
        RECT 0.090 729.980 689.780 732.180 ;
        RECT 0.090 728.820 0.700 729.980 ;
        RECT 4.300 728.820 689.780 729.980 ;
        RECT 0.090 726.620 689.780 728.820 ;
        RECT 0.090 725.460 685.700 726.620 ;
        RECT 689.300 725.460 689.780 726.620 ;
        RECT 0.090 723.260 689.780 725.460 ;
        RECT 0.090 722.100 0.700 723.260 ;
        RECT 4.300 722.100 689.780 723.260 ;
        RECT 0.090 719.900 689.780 722.100 ;
        RECT 0.090 718.740 685.700 719.900 ;
        RECT 689.300 718.740 689.780 719.900 ;
        RECT 0.090 716.540 689.780 718.740 ;
        RECT 0.090 715.380 0.700 716.540 ;
        RECT 4.300 715.380 689.780 716.540 ;
        RECT 0.090 713.180 689.780 715.380 ;
        RECT 0.090 712.020 685.700 713.180 ;
        RECT 689.300 712.020 689.780 713.180 ;
        RECT 0.090 709.820 689.780 712.020 ;
        RECT 0.090 708.660 0.700 709.820 ;
        RECT 4.300 708.660 689.780 709.820 ;
        RECT 0.090 706.460 689.780 708.660 ;
        RECT 0.090 705.300 685.700 706.460 ;
        RECT 689.300 705.300 689.780 706.460 ;
        RECT 0.090 703.100 689.780 705.300 ;
        RECT 0.090 701.940 0.700 703.100 ;
        RECT 4.300 701.940 689.780 703.100 ;
        RECT 0.090 699.740 689.780 701.940 ;
        RECT 0.090 698.580 685.700 699.740 ;
        RECT 689.300 698.580 689.780 699.740 ;
        RECT 0.090 696.380 689.780 698.580 ;
        RECT 0.090 695.220 0.700 696.380 ;
        RECT 4.300 695.220 689.780 696.380 ;
        RECT 0.090 689.660 689.780 695.220 ;
        RECT 0.090 688.500 685.700 689.660 ;
        RECT 689.300 688.500 689.780 689.660 ;
        RECT 0.090 686.300 689.780 688.500 ;
        RECT 0.090 685.140 0.700 686.300 ;
        RECT 4.300 685.140 689.780 686.300 ;
        RECT 0.090 682.940 689.780 685.140 ;
        RECT 0.090 681.780 685.700 682.940 ;
        RECT 689.300 681.780 689.780 682.940 ;
        RECT 0.090 679.580 689.780 681.780 ;
        RECT 0.090 678.420 0.700 679.580 ;
        RECT 4.300 678.420 689.780 679.580 ;
        RECT 0.090 676.220 689.780 678.420 ;
        RECT 0.090 675.060 685.700 676.220 ;
        RECT 689.300 675.060 689.780 676.220 ;
        RECT 0.090 672.860 689.780 675.060 ;
        RECT 0.090 671.700 0.700 672.860 ;
        RECT 4.300 671.700 689.780 672.860 ;
        RECT 0.090 669.500 689.780 671.700 ;
        RECT 0.090 668.340 685.700 669.500 ;
        RECT 689.300 668.340 689.780 669.500 ;
        RECT 0.090 666.140 689.780 668.340 ;
        RECT 0.090 664.980 0.700 666.140 ;
        RECT 4.300 664.980 689.780 666.140 ;
        RECT 0.090 662.780 689.780 664.980 ;
        RECT 0.090 661.620 685.700 662.780 ;
        RECT 689.300 661.620 689.780 662.780 ;
        RECT 0.090 659.420 689.780 661.620 ;
        RECT 0.090 658.260 0.700 659.420 ;
        RECT 4.300 658.260 689.780 659.420 ;
        RECT 0.090 656.060 689.780 658.260 ;
        RECT 0.090 654.900 685.700 656.060 ;
        RECT 689.300 654.900 689.780 656.060 ;
        RECT 0.090 652.700 689.780 654.900 ;
        RECT 0.090 651.540 0.700 652.700 ;
        RECT 4.300 651.540 689.780 652.700 ;
        RECT 0.090 649.340 689.780 651.540 ;
        RECT 0.090 648.180 685.700 649.340 ;
        RECT 689.300 648.180 689.780 649.340 ;
        RECT 0.090 645.980 689.780 648.180 ;
        RECT 0.090 644.820 0.700 645.980 ;
        RECT 4.300 644.820 689.780 645.980 ;
        RECT 0.090 642.620 689.780 644.820 ;
        RECT 0.090 641.460 685.700 642.620 ;
        RECT 689.300 641.460 689.780 642.620 ;
        RECT 0.090 635.900 689.780 641.460 ;
        RECT 0.090 634.740 0.700 635.900 ;
        RECT 4.300 634.740 689.780 635.900 ;
        RECT 0.090 632.540 689.780 634.740 ;
        RECT 0.090 631.380 685.700 632.540 ;
        RECT 689.300 631.380 689.780 632.540 ;
        RECT 0.090 629.180 689.780 631.380 ;
        RECT 0.090 628.020 0.700 629.180 ;
        RECT 4.300 628.020 689.780 629.180 ;
        RECT 0.090 625.820 689.780 628.020 ;
        RECT 0.090 624.660 685.700 625.820 ;
        RECT 689.300 624.660 689.780 625.820 ;
        RECT 0.090 622.460 689.780 624.660 ;
        RECT 0.090 621.300 0.700 622.460 ;
        RECT 4.300 621.300 689.780 622.460 ;
        RECT 0.090 619.100 689.780 621.300 ;
        RECT 0.090 617.940 685.700 619.100 ;
        RECT 689.300 617.940 689.780 619.100 ;
        RECT 0.090 615.740 689.780 617.940 ;
        RECT 0.090 614.580 0.700 615.740 ;
        RECT 4.300 614.580 689.780 615.740 ;
        RECT 0.090 612.380 689.780 614.580 ;
        RECT 0.090 611.220 685.700 612.380 ;
        RECT 689.300 611.220 689.780 612.380 ;
        RECT 0.090 609.020 689.780 611.220 ;
        RECT 0.090 607.860 0.700 609.020 ;
        RECT 4.300 607.860 689.780 609.020 ;
        RECT 0.090 605.660 689.780 607.860 ;
        RECT 0.090 604.500 685.700 605.660 ;
        RECT 689.300 604.500 689.780 605.660 ;
        RECT 0.090 602.300 689.780 604.500 ;
        RECT 0.090 601.140 0.700 602.300 ;
        RECT 4.300 601.140 689.780 602.300 ;
        RECT 0.090 598.940 689.780 601.140 ;
        RECT 0.090 597.780 685.700 598.940 ;
        RECT 689.300 597.780 689.780 598.940 ;
        RECT 0.090 595.580 689.780 597.780 ;
        RECT 0.090 594.420 0.700 595.580 ;
        RECT 4.300 594.420 689.780 595.580 ;
        RECT 0.090 592.220 689.780 594.420 ;
        RECT 0.090 591.060 685.700 592.220 ;
        RECT 689.300 591.060 689.780 592.220 ;
        RECT 0.090 588.860 689.780 591.060 ;
        RECT 0.090 587.700 0.700 588.860 ;
        RECT 4.300 587.700 689.780 588.860 ;
        RECT 0.090 582.140 689.780 587.700 ;
        RECT 0.090 580.980 685.700 582.140 ;
        RECT 689.300 580.980 689.780 582.140 ;
        RECT 0.090 578.780 689.780 580.980 ;
        RECT 0.090 577.620 0.700 578.780 ;
        RECT 4.300 577.620 689.780 578.780 ;
        RECT 0.090 575.420 689.780 577.620 ;
        RECT 0.090 574.260 685.700 575.420 ;
        RECT 689.300 574.260 689.780 575.420 ;
        RECT 0.090 572.060 689.780 574.260 ;
        RECT 0.090 570.900 0.700 572.060 ;
        RECT 4.300 570.900 689.780 572.060 ;
        RECT 0.090 568.700 689.780 570.900 ;
        RECT 0.090 567.540 685.700 568.700 ;
        RECT 689.300 567.540 689.780 568.700 ;
        RECT 0.090 565.340 689.780 567.540 ;
        RECT 0.090 564.180 0.700 565.340 ;
        RECT 4.300 564.180 689.780 565.340 ;
        RECT 0.090 561.980 689.780 564.180 ;
        RECT 0.090 560.820 685.700 561.980 ;
        RECT 689.300 560.820 689.780 561.980 ;
        RECT 0.090 558.620 689.780 560.820 ;
        RECT 0.090 557.460 0.700 558.620 ;
        RECT 4.300 557.460 689.780 558.620 ;
        RECT 0.090 555.260 689.780 557.460 ;
        RECT 0.090 554.100 685.700 555.260 ;
        RECT 689.300 554.100 689.780 555.260 ;
        RECT 0.090 551.900 689.780 554.100 ;
        RECT 0.090 550.740 0.700 551.900 ;
        RECT 4.300 550.740 689.780 551.900 ;
        RECT 0.090 548.540 689.780 550.740 ;
        RECT 0.090 547.380 685.700 548.540 ;
        RECT 689.300 547.380 689.780 548.540 ;
        RECT 0.090 545.180 689.780 547.380 ;
        RECT 0.090 544.020 0.700 545.180 ;
        RECT 4.300 544.020 689.780 545.180 ;
        RECT 0.090 541.820 689.780 544.020 ;
        RECT 0.090 540.660 685.700 541.820 ;
        RECT 689.300 540.660 689.780 541.820 ;
        RECT 0.090 538.460 689.780 540.660 ;
        RECT 0.090 537.300 0.700 538.460 ;
        RECT 4.300 537.300 689.780 538.460 ;
        RECT 0.090 535.100 689.780 537.300 ;
        RECT 0.090 533.940 685.700 535.100 ;
        RECT 689.300 533.940 689.780 535.100 ;
        RECT 0.090 528.380 689.780 533.940 ;
        RECT 0.090 527.220 0.700 528.380 ;
        RECT 4.300 527.220 689.780 528.380 ;
        RECT 0.090 525.020 689.780 527.220 ;
        RECT 0.090 523.860 685.700 525.020 ;
        RECT 689.300 523.860 689.780 525.020 ;
        RECT 0.090 521.660 689.780 523.860 ;
        RECT 0.090 520.500 0.700 521.660 ;
        RECT 4.300 520.500 689.780 521.660 ;
        RECT 0.090 518.300 689.780 520.500 ;
        RECT 0.090 517.140 685.700 518.300 ;
        RECT 689.300 517.140 689.780 518.300 ;
        RECT 0.090 514.940 689.780 517.140 ;
        RECT 0.090 513.780 0.700 514.940 ;
        RECT 4.300 513.780 689.780 514.940 ;
        RECT 0.090 511.580 689.780 513.780 ;
        RECT 0.090 510.420 685.700 511.580 ;
        RECT 689.300 510.420 689.780 511.580 ;
        RECT 0.090 508.220 689.780 510.420 ;
        RECT 0.090 507.060 0.700 508.220 ;
        RECT 4.300 507.060 689.780 508.220 ;
        RECT 0.090 504.860 689.780 507.060 ;
        RECT 0.090 503.700 685.700 504.860 ;
        RECT 689.300 503.700 689.780 504.860 ;
        RECT 0.090 501.500 689.780 503.700 ;
        RECT 0.090 500.340 0.700 501.500 ;
        RECT 4.300 500.340 689.780 501.500 ;
        RECT 0.090 498.140 689.780 500.340 ;
        RECT 0.090 496.980 685.700 498.140 ;
        RECT 689.300 496.980 689.780 498.140 ;
        RECT 0.090 494.780 689.780 496.980 ;
        RECT 0.090 493.620 0.700 494.780 ;
        RECT 4.300 493.620 689.780 494.780 ;
        RECT 0.090 491.420 689.780 493.620 ;
        RECT 0.090 490.260 685.700 491.420 ;
        RECT 689.300 490.260 689.780 491.420 ;
        RECT 0.090 488.060 689.780 490.260 ;
        RECT 0.090 486.900 0.700 488.060 ;
        RECT 4.300 486.900 689.780 488.060 ;
        RECT 0.090 484.700 689.780 486.900 ;
        RECT 0.090 483.540 685.700 484.700 ;
        RECT 689.300 483.540 689.780 484.700 ;
        RECT 0.090 481.340 689.780 483.540 ;
        RECT 0.090 480.180 0.700 481.340 ;
        RECT 4.300 480.180 689.780 481.340 ;
        RECT 0.090 474.620 689.780 480.180 ;
        RECT 0.090 473.460 685.700 474.620 ;
        RECT 689.300 473.460 689.780 474.620 ;
        RECT 0.090 471.260 689.780 473.460 ;
        RECT 0.090 470.100 0.700 471.260 ;
        RECT 4.300 470.100 689.780 471.260 ;
        RECT 0.090 467.900 689.780 470.100 ;
        RECT 0.090 466.740 685.700 467.900 ;
        RECT 689.300 466.740 689.780 467.900 ;
        RECT 0.090 464.540 689.780 466.740 ;
        RECT 0.090 463.380 0.700 464.540 ;
        RECT 4.300 463.380 689.780 464.540 ;
        RECT 0.090 461.180 689.780 463.380 ;
        RECT 0.090 460.020 685.700 461.180 ;
        RECT 689.300 460.020 689.780 461.180 ;
        RECT 0.090 457.820 689.780 460.020 ;
        RECT 0.090 456.660 0.700 457.820 ;
        RECT 4.300 456.660 689.780 457.820 ;
        RECT 0.090 454.460 689.780 456.660 ;
        RECT 0.090 453.300 685.700 454.460 ;
        RECT 689.300 453.300 689.780 454.460 ;
        RECT 0.090 451.100 689.780 453.300 ;
        RECT 0.090 449.940 0.700 451.100 ;
        RECT 4.300 449.940 689.780 451.100 ;
        RECT 0.090 447.740 689.780 449.940 ;
        RECT 0.090 446.580 685.700 447.740 ;
        RECT 689.300 446.580 689.780 447.740 ;
        RECT 0.090 444.380 689.780 446.580 ;
        RECT 0.090 443.220 0.700 444.380 ;
        RECT 4.300 443.220 689.780 444.380 ;
        RECT 0.090 441.020 689.780 443.220 ;
        RECT 0.090 439.860 685.700 441.020 ;
        RECT 689.300 439.860 689.780 441.020 ;
        RECT 0.090 437.660 689.780 439.860 ;
        RECT 0.090 436.500 0.700 437.660 ;
        RECT 4.300 436.500 689.780 437.660 ;
        RECT 0.090 434.300 689.780 436.500 ;
        RECT 0.090 433.140 685.700 434.300 ;
        RECT 689.300 433.140 689.780 434.300 ;
        RECT 0.090 430.940 689.780 433.140 ;
        RECT 0.090 429.780 0.700 430.940 ;
        RECT 4.300 429.780 689.780 430.940 ;
        RECT 0.090 427.580 689.780 429.780 ;
        RECT 0.090 426.420 685.700 427.580 ;
        RECT 689.300 426.420 689.780 427.580 ;
        RECT 0.090 420.860 689.780 426.420 ;
        RECT 0.090 419.700 0.700 420.860 ;
        RECT 4.300 419.700 689.780 420.860 ;
        RECT 0.090 417.500 689.780 419.700 ;
        RECT 0.090 416.340 685.700 417.500 ;
        RECT 689.300 416.340 689.780 417.500 ;
        RECT 0.090 414.140 689.780 416.340 ;
        RECT 0.090 412.980 0.700 414.140 ;
        RECT 4.300 412.980 689.780 414.140 ;
        RECT 0.090 410.780 689.780 412.980 ;
        RECT 0.090 409.620 685.700 410.780 ;
        RECT 689.300 409.620 689.780 410.780 ;
        RECT 0.090 407.420 689.780 409.620 ;
        RECT 0.090 406.260 0.700 407.420 ;
        RECT 4.300 406.260 689.780 407.420 ;
        RECT 0.090 404.060 689.780 406.260 ;
        RECT 0.090 402.900 685.700 404.060 ;
        RECT 689.300 402.900 689.780 404.060 ;
        RECT 0.090 400.700 689.780 402.900 ;
        RECT 0.090 399.540 0.700 400.700 ;
        RECT 4.300 399.540 689.780 400.700 ;
        RECT 0.090 397.340 689.780 399.540 ;
        RECT 0.090 396.180 685.700 397.340 ;
        RECT 689.300 396.180 689.780 397.340 ;
        RECT 0.090 393.980 689.780 396.180 ;
        RECT 0.090 392.820 0.700 393.980 ;
        RECT 4.300 392.820 689.780 393.980 ;
        RECT 0.090 390.620 689.780 392.820 ;
        RECT 0.090 389.460 685.700 390.620 ;
        RECT 689.300 389.460 689.780 390.620 ;
        RECT 0.090 387.260 689.780 389.460 ;
        RECT 0.090 386.100 0.700 387.260 ;
        RECT 4.300 386.100 689.780 387.260 ;
        RECT 0.090 383.900 689.780 386.100 ;
        RECT 0.090 382.740 685.700 383.900 ;
        RECT 689.300 382.740 689.780 383.900 ;
        RECT 0.090 380.540 689.780 382.740 ;
        RECT 0.090 379.380 0.700 380.540 ;
        RECT 4.300 379.380 689.780 380.540 ;
        RECT 0.090 377.180 689.780 379.380 ;
        RECT 0.090 376.020 685.700 377.180 ;
        RECT 689.300 376.020 689.780 377.180 ;
        RECT 0.090 370.460 689.780 376.020 ;
        RECT 0.090 369.300 0.700 370.460 ;
        RECT 4.300 369.300 689.780 370.460 ;
        RECT 0.090 367.100 689.780 369.300 ;
        RECT 0.090 365.940 685.700 367.100 ;
        RECT 689.300 365.940 689.780 367.100 ;
        RECT 0.090 363.740 689.780 365.940 ;
        RECT 0.090 362.580 0.700 363.740 ;
        RECT 4.300 362.580 689.780 363.740 ;
        RECT 0.090 360.380 689.780 362.580 ;
        RECT 0.090 359.220 685.700 360.380 ;
        RECT 689.300 359.220 689.780 360.380 ;
        RECT 0.090 357.020 689.780 359.220 ;
        RECT 0.090 355.860 0.700 357.020 ;
        RECT 4.300 355.860 689.780 357.020 ;
        RECT 0.090 353.660 689.780 355.860 ;
        RECT 0.090 352.500 685.700 353.660 ;
        RECT 689.300 352.500 689.780 353.660 ;
        RECT 0.090 350.300 689.780 352.500 ;
        RECT 0.090 349.140 0.700 350.300 ;
        RECT 4.300 349.140 689.780 350.300 ;
        RECT 0.090 346.940 689.780 349.140 ;
        RECT 0.090 345.780 685.700 346.940 ;
        RECT 689.300 345.780 689.780 346.940 ;
        RECT 0.090 343.580 689.780 345.780 ;
        RECT 0.090 342.420 0.700 343.580 ;
        RECT 4.300 342.420 689.780 343.580 ;
        RECT 0.090 340.220 689.780 342.420 ;
        RECT 0.090 339.060 685.700 340.220 ;
        RECT 689.300 339.060 689.780 340.220 ;
        RECT 0.090 336.860 689.780 339.060 ;
        RECT 0.090 335.700 0.700 336.860 ;
        RECT 4.300 335.700 689.780 336.860 ;
        RECT 0.090 333.500 689.780 335.700 ;
        RECT 0.090 332.340 685.700 333.500 ;
        RECT 689.300 332.340 689.780 333.500 ;
        RECT 0.090 330.140 689.780 332.340 ;
        RECT 0.090 328.980 0.700 330.140 ;
        RECT 4.300 328.980 689.780 330.140 ;
        RECT 0.090 326.780 689.780 328.980 ;
        RECT 0.090 325.620 685.700 326.780 ;
        RECT 689.300 325.620 689.780 326.780 ;
        RECT 0.090 323.420 689.780 325.620 ;
        RECT 0.090 322.260 0.700 323.420 ;
        RECT 4.300 322.260 689.780 323.420 ;
        RECT 0.090 316.700 689.780 322.260 ;
        RECT 0.090 315.540 685.700 316.700 ;
        RECT 689.300 315.540 689.780 316.700 ;
        RECT 0.090 313.340 689.780 315.540 ;
        RECT 0.090 312.180 0.700 313.340 ;
        RECT 4.300 312.180 689.780 313.340 ;
        RECT 0.090 309.980 689.780 312.180 ;
        RECT 0.090 308.820 685.700 309.980 ;
        RECT 689.300 308.820 689.780 309.980 ;
        RECT 0.090 306.620 689.780 308.820 ;
        RECT 0.090 305.460 0.700 306.620 ;
        RECT 4.300 305.460 689.780 306.620 ;
        RECT 0.090 303.260 689.780 305.460 ;
        RECT 0.090 302.100 685.700 303.260 ;
        RECT 689.300 302.100 689.780 303.260 ;
        RECT 0.090 299.900 689.780 302.100 ;
        RECT 0.090 298.740 0.700 299.900 ;
        RECT 4.300 298.740 689.780 299.900 ;
        RECT 0.090 296.540 689.780 298.740 ;
        RECT 0.090 295.380 685.700 296.540 ;
        RECT 689.300 295.380 689.780 296.540 ;
        RECT 0.090 293.180 689.780 295.380 ;
        RECT 0.090 292.020 0.700 293.180 ;
        RECT 4.300 292.020 689.780 293.180 ;
        RECT 0.090 289.820 689.780 292.020 ;
        RECT 0.090 288.660 685.700 289.820 ;
        RECT 689.300 288.660 689.780 289.820 ;
        RECT 0.090 286.460 689.780 288.660 ;
        RECT 0.090 285.300 0.700 286.460 ;
        RECT 4.300 285.300 689.780 286.460 ;
        RECT 0.090 283.100 689.780 285.300 ;
        RECT 0.090 281.940 685.700 283.100 ;
        RECT 689.300 281.940 689.780 283.100 ;
        RECT 0.090 279.740 689.780 281.940 ;
        RECT 0.090 278.580 0.700 279.740 ;
        RECT 4.300 278.580 689.780 279.740 ;
        RECT 0.090 276.380 689.780 278.580 ;
        RECT 0.090 275.220 685.700 276.380 ;
        RECT 689.300 275.220 689.780 276.380 ;
        RECT 0.090 273.020 689.780 275.220 ;
        RECT 0.090 271.860 0.700 273.020 ;
        RECT 4.300 271.860 689.780 273.020 ;
        RECT 0.090 269.660 689.780 271.860 ;
        RECT 0.090 268.500 685.700 269.660 ;
        RECT 689.300 268.500 689.780 269.660 ;
        RECT 0.090 262.940 689.780 268.500 ;
        RECT 0.090 261.780 0.700 262.940 ;
        RECT 4.300 261.780 689.780 262.940 ;
        RECT 0.090 259.580 689.780 261.780 ;
        RECT 0.090 258.420 685.700 259.580 ;
        RECT 689.300 258.420 689.780 259.580 ;
        RECT 0.090 256.220 689.780 258.420 ;
        RECT 0.090 255.060 0.700 256.220 ;
        RECT 4.300 255.060 689.780 256.220 ;
        RECT 0.090 252.860 689.780 255.060 ;
        RECT 0.090 251.700 685.700 252.860 ;
        RECT 689.300 251.700 689.780 252.860 ;
        RECT 0.090 249.500 689.780 251.700 ;
        RECT 0.090 248.340 0.700 249.500 ;
        RECT 4.300 248.340 689.780 249.500 ;
        RECT 0.090 246.140 689.780 248.340 ;
        RECT 0.090 244.980 685.700 246.140 ;
        RECT 689.300 244.980 689.780 246.140 ;
        RECT 0.090 242.780 689.780 244.980 ;
        RECT 0.090 241.620 0.700 242.780 ;
        RECT 4.300 241.620 689.780 242.780 ;
        RECT 0.090 239.420 689.780 241.620 ;
        RECT 0.090 238.260 685.700 239.420 ;
        RECT 689.300 238.260 689.780 239.420 ;
        RECT 0.090 236.060 689.780 238.260 ;
        RECT 0.090 234.900 0.700 236.060 ;
        RECT 4.300 234.900 689.780 236.060 ;
        RECT 0.090 232.700 689.780 234.900 ;
        RECT 0.090 231.540 685.700 232.700 ;
        RECT 689.300 231.540 689.780 232.700 ;
        RECT 0.090 229.340 689.780 231.540 ;
        RECT 0.090 228.180 0.700 229.340 ;
        RECT 4.300 228.180 689.780 229.340 ;
        RECT 0.090 225.980 689.780 228.180 ;
        RECT 0.090 224.820 685.700 225.980 ;
        RECT 689.300 224.820 689.780 225.980 ;
        RECT 0.090 222.620 689.780 224.820 ;
        RECT 0.090 221.460 0.700 222.620 ;
        RECT 4.300 221.460 689.780 222.620 ;
        RECT 0.090 219.260 689.780 221.460 ;
        RECT 0.090 218.100 685.700 219.260 ;
        RECT 689.300 218.100 689.780 219.260 ;
        RECT 0.090 215.900 689.780 218.100 ;
        RECT 0.090 214.740 0.700 215.900 ;
        RECT 4.300 214.740 689.780 215.900 ;
        RECT 0.090 209.180 689.780 214.740 ;
        RECT 0.090 208.020 685.700 209.180 ;
        RECT 689.300 208.020 689.780 209.180 ;
        RECT 0.090 205.820 689.780 208.020 ;
        RECT 0.090 204.660 0.700 205.820 ;
        RECT 4.300 204.660 689.780 205.820 ;
        RECT 0.090 202.460 689.780 204.660 ;
        RECT 0.090 201.300 685.700 202.460 ;
        RECT 689.300 201.300 689.780 202.460 ;
        RECT 0.090 199.100 689.780 201.300 ;
        RECT 0.090 197.940 0.700 199.100 ;
        RECT 4.300 197.940 689.780 199.100 ;
        RECT 0.090 195.740 689.780 197.940 ;
        RECT 0.090 194.580 685.700 195.740 ;
        RECT 689.300 194.580 689.780 195.740 ;
        RECT 0.090 192.380 689.780 194.580 ;
        RECT 0.090 191.220 0.700 192.380 ;
        RECT 4.300 191.220 689.780 192.380 ;
        RECT 0.090 189.020 689.780 191.220 ;
        RECT 0.090 187.860 685.700 189.020 ;
        RECT 689.300 187.860 689.780 189.020 ;
        RECT 0.090 185.660 689.780 187.860 ;
        RECT 0.090 184.500 0.700 185.660 ;
        RECT 4.300 184.500 689.780 185.660 ;
        RECT 0.090 182.300 689.780 184.500 ;
        RECT 0.090 181.140 685.700 182.300 ;
        RECT 689.300 181.140 689.780 182.300 ;
        RECT 0.090 178.940 689.780 181.140 ;
        RECT 0.090 177.780 0.700 178.940 ;
        RECT 4.300 177.780 689.780 178.940 ;
        RECT 0.090 175.580 689.780 177.780 ;
        RECT 0.090 174.420 685.700 175.580 ;
        RECT 689.300 174.420 689.780 175.580 ;
        RECT 0.090 172.220 689.780 174.420 ;
        RECT 0.090 171.060 0.700 172.220 ;
        RECT 4.300 171.060 689.780 172.220 ;
        RECT 0.090 168.860 689.780 171.060 ;
        RECT 0.090 167.700 685.700 168.860 ;
        RECT 689.300 167.700 689.780 168.860 ;
        RECT 0.090 165.500 689.780 167.700 ;
        RECT 0.090 164.340 0.700 165.500 ;
        RECT 4.300 164.340 689.780 165.500 ;
        RECT 0.090 162.140 689.780 164.340 ;
        RECT 0.090 160.980 685.700 162.140 ;
        RECT 689.300 160.980 689.780 162.140 ;
        RECT 0.090 155.420 689.780 160.980 ;
        RECT 0.090 154.260 0.700 155.420 ;
        RECT 4.300 154.260 689.780 155.420 ;
        RECT 0.090 152.060 689.780 154.260 ;
        RECT 0.090 150.900 685.700 152.060 ;
        RECT 689.300 150.900 689.780 152.060 ;
        RECT 0.090 148.700 689.780 150.900 ;
        RECT 0.090 147.540 0.700 148.700 ;
        RECT 4.300 147.540 689.780 148.700 ;
        RECT 0.090 145.340 689.780 147.540 ;
        RECT 0.090 144.180 685.700 145.340 ;
        RECT 689.300 144.180 689.780 145.340 ;
        RECT 0.090 141.980 689.780 144.180 ;
        RECT 0.090 140.820 0.700 141.980 ;
        RECT 4.300 140.820 689.780 141.980 ;
        RECT 0.090 138.620 689.780 140.820 ;
        RECT 0.090 137.460 685.700 138.620 ;
        RECT 689.300 137.460 689.780 138.620 ;
        RECT 0.090 135.260 689.780 137.460 ;
        RECT 0.090 134.100 0.700 135.260 ;
        RECT 4.300 134.100 689.780 135.260 ;
        RECT 0.090 131.900 689.780 134.100 ;
        RECT 0.090 130.740 685.700 131.900 ;
        RECT 689.300 130.740 689.780 131.900 ;
        RECT 0.090 128.540 689.780 130.740 ;
        RECT 0.090 127.380 0.700 128.540 ;
        RECT 4.300 127.380 689.780 128.540 ;
        RECT 0.090 125.180 689.780 127.380 ;
        RECT 0.090 124.020 685.700 125.180 ;
        RECT 689.300 124.020 689.780 125.180 ;
        RECT 0.090 121.820 689.780 124.020 ;
        RECT 0.090 120.660 0.700 121.820 ;
        RECT 4.300 120.660 689.780 121.820 ;
        RECT 0.090 118.460 689.780 120.660 ;
        RECT 0.090 117.300 685.700 118.460 ;
        RECT 689.300 117.300 689.780 118.460 ;
        RECT 0.090 115.100 689.780 117.300 ;
        RECT 0.090 113.940 0.700 115.100 ;
        RECT 4.300 113.940 689.780 115.100 ;
        RECT 0.090 111.740 689.780 113.940 ;
        RECT 0.090 110.580 685.700 111.740 ;
        RECT 689.300 110.580 689.780 111.740 ;
        RECT 0.090 108.380 689.780 110.580 ;
        RECT 0.090 107.220 0.700 108.380 ;
        RECT 4.300 107.220 689.780 108.380 ;
        RECT 0.090 101.660 689.780 107.220 ;
        RECT 0.090 100.500 685.700 101.660 ;
        RECT 689.300 100.500 689.780 101.660 ;
        RECT 0.090 98.300 689.780 100.500 ;
        RECT 0.090 97.140 0.700 98.300 ;
        RECT 4.300 97.140 689.780 98.300 ;
        RECT 0.090 94.940 689.780 97.140 ;
        RECT 0.090 93.780 685.700 94.940 ;
        RECT 689.300 93.780 689.780 94.940 ;
        RECT 0.090 91.580 689.780 93.780 ;
        RECT 0.090 90.420 0.700 91.580 ;
        RECT 4.300 90.420 689.780 91.580 ;
        RECT 0.090 88.220 689.780 90.420 ;
        RECT 0.090 87.060 685.700 88.220 ;
        RECT 689.300 87.060 689.780 88.220 ;
        RECT 0.090 84.860 689.780 87.060 ;
        RECT 0.090 83.700 0.700 84.860 ;
        RECT 4.300 83.700 689.780 84.860 ;
        RECT 0.090 81.500 689.780 83.700 ;
        RECT 0.090 80.340 685.700 81.500 ;
        RECT 689.300 80.340 689.780 81.500 ;
        RECT 0.090 78.140 689.780 80.340 ;
        RECT 0.090 76.980 0.700 78.140 ;
        RECT 4.300 76.980 689.780 78.140 ;
        RECT 0.090 74.780 689.780 76.980 ;
        RECT 0.090 73.620 685.700 74.780 ;
        RECT 689.300 73.620 689.780 74.780 ;
        RECT 0.090 71.420 689.780 73.620 ;
        RECT 0.090 70.260 0.700 71.420 ;
        RECT 4.300 70.260 689.780 71.420 ;
        RECT 0.090 68.060 689.780 70.260 ;
        RECT 0.090 66.900 685.700 68.060 ;
        RECT 689.300 66.900 689.780 68.060 ;
        RECT 0.090 64.700 689.780 66.900 ;
        RECT 0.090 63.540 0.700 64.700 ;
        RECT 4.300 63.540 689.780 64.700 ;
        RECT 0.090 61.340 689.780 63.540 ;
        RECT 0.090 60.180 685.700 61.340 ;
        RECT 689.300 60.180 689.780 61.340 ;
        RECT 0.090 57.980 689.780 60.180 ;
        RECT 0.090 56.820 0.700 57.980 ;
        RECT 4.300 56.820 689.780 57.980 ;
        RECT 0.090 54.620 689.780 56.820 ;
        RECT 0.090 53.460 685.700 54.620 ;
        RECT 689.300 53.460 689.780 54.620 ;
        RECT 0.090 47.900 689.780 53.460 ;
        RECT 0.090 46.740 0.700 47.900 ;
        RECT 4.300 46.740 689.780 47.900 ;
        RECT 0.090 44.540 689.780 46.740 ;
        RECT 0.090 43.380 685.700 44.540 ;
        RECT 689.300 43.380 689.780 44.540 ;
        RECT 0.090 41.180 689.780 43.380 ;
        RECT 0.090 40.020 0.700 41.180 ;
        RECT 4.300 40.020 689.780 41.180 ;
        RECT 0.090 37.820 689.780 40.020 ;
        RECT 0.090 36.660 685.700 37.820 ;
        RECT 689.300 36.660 689.780 37.820 ;
        RECT 0.090 34.460 689.780 36.660 ;
        RECT 0.090 33.300 0.700 34.460 ;
        RECT 4.300 33.300 689.780 34.460 ;
        RECT 0.090 31.100 689.780 33.300 ;
        RECT 0.090 29.940 685.700 31.100 ;
        RECT 689.300 29.940 689.780 31.100 ;
        RECT 0.090 27.740 689.780 29.940 ;
        RECT 0.090 26.580 0.700 27.740 ;
        RECT 4.300 26.580 689.780 27.740 ;
        RECT 0.090 24.380 689.780 26.580 ;
        RECT 0.090 23.220 685.700 24.380 ;
        RECT 689.300 23.220 689.780 24.380 ;
        RECT 0.090 21.020 689.780 23.220 ;
        RECT 0.090 19.860 0.700 21.020 ;
        RECT 4.300 19.860 689.780 21.020 ;
        RECT 0.090 17.660 689.780 19.860 ;
        RECT 0.090 16.500 685.700 17.660 ;
        RECT 689.300 16.500 689.780 17.660 ;
        RECT 0.090 14.300 689.780 16.500 ;
        RECT 0.090 13.140 0.700 14.300 ;
        RECT 4.300 13.140 689.780 14.300 ;
        RECT 0.090 10.940 689.780 13.140 ;
        RECT 0.090 9.780 685.700 10.940 ;
        RECT 689.300 9.780 689.780 10.940 ;
        RECT 0.090 7.580 689.780 9.780 ;
        RECT 0.090 6.420 0.700 7.580 ;
        RECT 4.300 6.420 689.780 7.580 ;
        RECT 0.090 4.220 689.780 6.420 ;
        RECT 0.090 3.500 685.700 4.220 ;
        RECT 689.300 3.500 689.780 4.220 ;
      LAYER Metal4 ;
        RECT 18.620 15.080 21.940 765.430 ;
        RECT 24.140 15.080 98.740 765.430 ;
        RECT 100.940 15.080 175.540 765.430 ;
        RECT 177.740 15.080 252.340 765.430 ;
        RECT 254.540 15.080 329.140 765.430 ;
        RECT 331.340 15.080 405.940 765.430 ;
        RECT 408.140 15.080 482.740 765.430 ;
        RECT 484.940 15.080 559.540 765.430 ;
        RECT 561.740 15.080 636.340 765.430 ;
        RECT 638.540 15.080 661.780 765.430 ;
        RECT 18.620 13.530 661.780 15.080 ;
  END
END tiny_user_project
END LIBRARY

