VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO serv_0
  CLASS BLOCK ;
  FOREIGN serv_0 ;
  ORIGIN 0.000 0.000 ;
  SIZE 700.000 BY 600.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 698.000 21.280 700.000 21.840 ;
    END
  END io_in[0]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 698.000 61.040 700.000 61.600 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 698.000 100.800 700.000 101.360 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 698.000 140.560 700.000 141.120 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 698.000 180.320 700.000 180.880 ;
    END
  END io_in[4]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 698.000 418.880 700.000 419.440 ;
    END
  END io_oeb[0]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 698.000 458.640 700.000 459.200 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 698.000 498.400 700.000 498.960 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 698.000 538.160 700.000 538.720 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 698.000 577.920 700.000 578.480 ;
    END
  END io_oeb[4]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 698.000 220.080 700.000 220.640 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 698.000 259.840 700.000 260.400 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 698.000 299.600 700.000 300.160 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 698.000 339.360 700.000 339.920 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 698.000 379.120 700.000 379.680 ;
    END
  END io_out[4]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 67.240 15.380 68.840 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 112.240 15.380 113.840 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 157.240 15.380 158.840 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 202.240 15.380 203.840 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 247.240 15.380 248.840 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 292.240 15.380 293.840 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 337.240 15.380 338.840 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 382.240 15.380 383.840 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 427.240 15.380 428.840 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 472.240 15.380 473.840 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 517.240 15.380 518.840 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 562.240 15.380 563.840 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 607.240 15.380 608.840 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 652.240 15.380 653.840 584.380 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 44.740 15.380 46.340 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 89.740 15.380 91.340 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 134.740 15.380 136.340 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 179.740 15.380 181.340 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 224.740 15.380 226.340 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 269.740 15.380 271.340 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 314.740 15.380 316.340 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 359.740 15.380 361.340 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 404.740 15.380 406.340 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 449.740 15.380 451.340 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 494.740 15.380 496.340 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 539.740 15.380 541.340 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 584.740 15.380 586.340 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 629.740 15.380 631.340 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 674.740 15.380 676.340 584.380 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 693.280 584.380 ;
      LAYER Metal2 ;
        RECT 22.380 3.450 698.740 584.270 ;
      LAYER Metal3 ;
        RECT 22.330 578.780 698.790 584.220 ;
        RECT 22.330 577.620 697.700 578.780 ;
        RECT 22.330 539.020 698.790 577.620 ;
        RECT 22.330 537.860 697.700 539.020 ;
        RECT 22.330 499.260 698.790 537.860 ;
        RECT 22.330 498.100 697.700 499.260 ;
        RECT 22.330 459.500 698.790 498.100 ;
        RECT 22.330 458.340 697.700 459.500 ;
        RECT 22.330 419.740 698.790 458.340 ;
        RECT 22.330 418.580 697.700 419.740 ;
        RECT 22.330 379.980 698.790 418.580 ;
        RECT 22.330 378.820 697.700 379.980 ;
        RECT 22.330 340.220 698.790 378.820 ;
        RECT 22.330 339.060 697.700 340.220 ;
        RECT 22.330 300.460 698.790 339.060 ;
        RECT 22.330 299.300 697.700 300.460 ;
        RECT 22.330 260.700 698.790 299.300 ;
        RECT 22.330 259.540 697.700 260.700 ;
        RECT 22.330 220.940 698.790 259.540 ;
        RECT 22.330 219.780 697.700 220.940 ;
        RECT 22.330 181.180 698.790 219.780 ;
        RECT 22.330 180.020 697.700 181.180 ;
        RECT 22.330 141.420 698.790 180.020 ;
        RECT 22.330 140.260 697.700 141.420 ;
        RECT 22.330 101.660 698.790 140.260 ;
        RECT 22.330 100.500 697.700 101.660 ;
        RECT 22.330 61.900 698.790 100.500 ;
        RECT 22.330 60.740 697.700 61.900 ;
        RECT 22.330 22.140 698.790 60.740 ;
        RECT 22.330 20.980 697.700 22.140 ;
        RECT 22.330 3.500 698.790 20.980 ;
      LAYER Metal4 ;
        RECT 429.660 15.080 449.440 496.070 ;
        RECT 451.640 15.080 471.940 496.070 ;
        RECT 474.140 15.080 494.440 496.070 ;
        RECT 496.640 15.080 516.940 496.070 ;
        RECT 519.140 15.080 539.440 496.070 ;
        RECT 541.640 15.080 561.940 496.070 ;
        RECT 564.140 15.080 584.440 496.070 ;
        RECT 586.640 15.080 606.940 496.070 ;
        RECT 609.140 15.080 629.440 496.070 ;
        RECT 631.640 15.080 651.940 496.070 ;
        RECT 654.140 15.080 674.440 496.070 ;
        RECT 676.640 15.080 688.660 496.070 ;
        RECT 429.660 3.450 688.660 15.080 ;
  END
END serv_0
END LIBRARY

